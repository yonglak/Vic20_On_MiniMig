-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity cart_rom is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of cart_rom is


  type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"0F",x"A0",x"09",x"A0",x"41",x"30",x"C3",x"C2", -- 0x0000 --41
    x"CD",x"68",x"A8",x"68",x"AA",x"68",x"40",x"78", -- 0x0008
    x"D8",x"A2",x"FF",x"9A",x"20",x"8A",x"FF",x"A9", -- 0x0010
    x"00",x"8D",x"1E",x"91",x"A9",x"C0",x"8D",x"2E", -- 0x0018
    x"91",x"A9",x"40",x"8D",x"1B",x"91",x"8D",x"2B", -- 0x0020
    x"91",x"A9",x"FF",x"8D",x"22",x"91",x"A9",x"80", -- 0x0028
    x"8D",x"13",x"91",x"D8",x"78",x"A9",x"00",x"8D", -- 0x0030
    x"1E",x"91",x"8D",x"2E",x"91",x"AD",x"1C",x"91", -- 0x0038
    x"29",x"3F",x"8D",x"1C",x"91",x"A9",x"80",x"85", -- 0x0040
    x"89",x"85",x"8A",x"85",x"8B",x"85",x"8C",x"A9", -- 0x0048
    x"00",x"85",x"8D",x"85",x"52",x"85",x"53",x"85", -- 0x0050
    x"51",x"A9",x"4C",x"85",x"59",x"A2",x"00",x"A9", -- 0x0058
    x"20",x"9D",x"00",x"1E",x"9D",x"00",x"1F",x"E8", -- 0x0060
    x"D0",x"F7",x"A2",x"0F",x"BD",x"AC",x"A0",x"9D", -- 0x0068
    x"00",x"90",x"CA",x"10",x"F7",x"E8",x"BD",x"00", -- 0x0070
    x"80",x"9D",x"00",x"10",x"BD",x"00",x"81",x"9D", -- 0x0078
    x"00",x"11",x"CA",x"D0",x"F1",x"20",x"9F",x"A4", -- 0x0080
    x"A2",x"10",x"BD",x"2A",x"BE",x"9D",x"00",x"1E", -- 0x0088
    x"CA",x"10",x"F7",x"A2",x"77",x"BD",x"3B",x"BE", -- 0x0090
    x"9D",x"78",x"14",x"CA",x"10",x"F7",x"20",x"CF", -- 0x0098
    x"A0",x"20",x"56",x"A2",x"A2",x"0C",x"20",x"F2", -- 0x00A0
    x"A4",x"4C",x"7C",x"A1",x"02",x"19",x"97",x"2C", -- 0x00A8
    x"00",x"FC",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00B0
    x"00",x"00",x"00",x"08",x"A9",x"00",x"A2",x"04", -- 0x00B8
    x"95",x"1D",x"CA",x"10",x"FB",x"A9",x"03",x"85", -- 0x00C0
    x"44",x"20",x"EA",x"B1",x"20",x"39",x"B1",x"A2", -- 0x00C8
    x"00",x"A9",x"00",x"85",x"2D",x"A4",x"2D",x"B9", -- 0x00D0
    x"9F",x"B4",x"85",x"2B",x"B9",x"A4",x"B4",x"85", -- 0x00D8
    x"2C",x"A9",x"0B",x"85",x"2E",x"BD",x"A9",x"B4", -- 0x00E0
    x"9D",x"78",x"18",x"A4",x"1D",x"A5",x"2C",x"18", -- 0x00E8
    x"79",x"E5",x"B4",x"9D",x"3C",x"18",x"A5",x"2B", -- 0x00F0
    x"9D",x"00",x"18",x"69",x"10",x"85",x"2B",x"E8", -- 0x00F8
    x"C6",x"2E",x"10",x"E1",x"E6",x"2D",x"E0",x"3C", -- 0x0100
    x"D0",x"CB",x"A2",x"00",x"A0",x"12",x"96",x"06", -- 0x0108
    x"88",x"10",x"FB",x"E8",x"A0",x"04",x"96",x"18", -- 0x0110
    x"88",x"10",x"FB",x"86",x"11",x"E8",x"86",x"4B", -- 0x0118
    x"A9",x"32",x"85",x"24",x"A9",x"03",x"85",x"2F", -- 0x0120
    x"A6",x"1D",x"BD",x"EE",x"B4",x"85",x"54",x"BD", -- 0x0128
    x"F7",x"B4",x"85",x"55",x"A2",x"09",x"BD",x"30", -- 0x0130
    x"B7",x"95",x"7F",x"CA",x"10",x"F8",x"20",x"2D", -- 0x0138
    x"A2",x"A2",x"3F",x"BD",x"6B",x"B7",x"9D",x"40", -- 0x0140
    x"13",x"9D",x"80",x"13",x"9D",x"C0",x"13",x"9D", -- 0x0148
    x"00",x"14",x"CA",x"10",x"EE",x"A0",x"1F",x"A9", -- 0x0150
    x"87",x"BE",x"AB",x"B7",x"9D",x"89",x"1F",x"38", -- 0x0158
    x"E9",x"01",x"88",x"10",x"F4",x"A9",x"09",x"85", -- 0x0160
    x"3F",x"A9",x"0B",x"85",x"40",x"A9",x"FA",x"85", -- 0x0168
    x"41",x"A2",x"0C",x"20",x"F2",x"A4",x"20",x"9F", -- 0x0170
    x"A4",x"4C",x"63",x"A4",x"A9",x"86",x"8D",x"14", -- 0x0178
    x"91",x"A9",x"42",x"8D",x"15",x"91",x"20",x"92", -- 0x0180
    x"A1",x"AD",x"1D",x"91",x"29",x"40",x"F0",x"F9", -- 0x0188
    x"D0",x"EA",x"A9",x"00",x"85",x"37",x"A6",x"37", -- 0x0190
    x"E6",x"09",x"B5",x"7F",x"30",x"18",x"F0",x"05", -- 0x0198
    x"D6",x"7F",x"4C",x"B6",x"A1",x"BD",x"5A",x"B7", -- 0x01A0
    x"C9",x"FF",x"F0",x"0E",x"85",x"5B",x"BD",x"4C", -- 0x01A8
    x"B7",x"85",x"5A",x"20",x"59",x"00",x"E6",x"37", -- 0x01B0
    x"D0",x"DC",x"A5",x"44",x"F0",x"33",x"A5",x"0B", -- 0x01B8
    x"F0",x"03",x"4C",x"D6",x"A3",x"A5",x"24",x"D0", -- 0x01C0
    x"27",x"20",x"81",x"A4",x"A5",x"14",x"05",x"15", -- 0x01C8
    x"05",x"16",x"05",x"17",x"05",x"81",x"D0",x"18", -- 0x01D0
    x"A5",x"87",x"10",x"14",x"E6",x"1D",x"A5",x"1D", -- 0x01D8
    x"C9",x"09",x"D0",x"02",x"A9",x"01",x"85",x"1D", -- 0x01E0
    x"A2",x"32",x"20",x"F2",x"A4",x"4C",x"CF",x"A0", -- 0x01E8
    x"60",x"A5",x"1F",x"F0",x"0A",x"A5",x"81",x"C9", -- 0x01F0
    x"14",x"D0",x"03",x"4C",x"56",x"A2",x"60",x"A5", -- 0x01F8
    x"89",x"10",x"29",x"A9",x"80",x"A2",x"09",x"95", -- 0x0200
    x"7F",x"CA",x"10",x"FB",x"A9",x"00",x"85",x"89", -- 0x0208
    x"85",x"2B",x"20",x"81",x"A4",x"A5",x"20",x"C5", -- 0x0210
    x"52",x"A5",x"21",x"E5",x"53",x"90",x"0D",x"A5", -- 0x0218
    x"20",x"85",x"52",x"A5",x"21",x"85",x"53",x"A2", -- 0x0220
    x"08",x"4C",x"49",x"B1",x"60",x"A2",x"00",x"A9", -- 0x0228
    x"20",x"9D",x"17",x"1E",x"9D",x"17",x"1F",x"CA", -- 0x0230
    x"D0",x"F7",x"60",x"A9",x"06",x"85",x"89",x"A6", -- 0x0238
    x"2B",x"E6",x"2B",x"E0",x"14",x"F0",x"0B",x"E0", -- 0x0240
    x"09",x"B0",x"06",x"BD",x"1B",x"BD",x"9D",x"1E", -- 0x0248
    x"1E",x"60",x"A9",x"80",x"85",x"89",x"A2",x"00", -- 0x0250
    x"86",x"8C",x"86",x"8A",x"86",x"44",x"86",x"11", -- 0x0258
    x"E8",x"86",x"1F",x"A9",x"80",x"A2",x"0A",x"95", -- 0x0260
    x"7F",x"CA",x"10",x"FB",x"85",x"8B",x"20",x"2D", -- 0x0268
    x"A2",x"A9",x"9D",x"A2",x"0E",x"9D",x"E7",x"1F", -- 0x0270
    x"38",x"E9",x"01",x"CA",x"10",x"F7",x"20",x"DF", -- 0x0278
    x"A4",x"A9",x"00",x"85",x"33",x"A9",x"0A",x"85", -- 0x0280
    x"34",x"A2",x"03",x"20",x"F2",x"A4",x"A2",x"07", -- 0x0288
    x"20",x"F2",x"A4",x"A2",x"0B",x"20",x"F2",x"A4", -- 0x0290
    x"A2",x"23",x"4C",x"F2",x"A4",x"A4",x"29",x"B9", -- 0x0298
    x"EE",x"B3",x"85",x"00",x"B9",x"07",x"B4",x"85", -- 0x02A0
    x"01",x"A6",x"33",x"E6",x"33",x"BD",x"24",x"BD", -- 0x02A8
    x"C9",x"C0",x"B0",x"0D",x"A4",x"28",x"91",x"00", -- 0x02B0
    x"E6",x"28",x"A5",x"34",x"F0",x"DF",x"85",x"8A", -- 0x02B8
    x"60",x"C9",x"FF",x"F0",x"1E",x"C9",x"FE",x"F0", -- 0x02C0
    x"12",x"BD",x"25",x"BD",x"85",x"28",x"BD",x"26", -- 0x02C8
    x"BD",x"85",x"29",x"E8",x"E8",x"E8",x"86",x"33", -- 0x02D0
    x"4C",x"9D",x"A2",x"BD",x"25",x"BD",x"85",x"34", -- 0x02D8
    x"E6",x"33",x"60",x"A2",x"00",x"86",x"1D",x"E8", -- 0x02E0
    x"86",x"48",x"86",x"49",x"86",x"4A",x"20",x"CF", -- 0x02E8
    x"A0",x"20",x"81",x"A4",x"A9",x"64",x"85",x"8B", -- 0x02F0
    x"A9",x"80",x"85",x"8A",x"85",x"84",x"A5",x"20", -- 0x02F8
    x"85",x"09",x"60",x"A5",x"87",x"30",x"01",x"60", -- 0x0300
    x"A5",x"17",x"D0",x"03",x"20",x"94",x"A7",x"C6", -- 0x0308
    x"48",x"D0",x"1B",x"E6",x"4E",x"A6",x"4E",x"BD", -- 0x0310
    x"16",x"BA",x"29",x"0F",x"85",x"48",x"BD",x"18", -- 0x0318
    x"BA",x"4A",x"90",x"06",x"A5",x"49",x"85",x"4A", -- 0x0320
    x"B0",x"04",x"A9",x"00",x"85",x"4A",x"A5",x"2F", -- 0x0328
    x"18",x"65",x"4A",x"C9",x"03",x"90",x"04",x"C9", -- 0x0330
    x"98",x"90",x"0C",x"A5",x"49",x"49",x"FF",x"18", -- 0x0338
    x"69",x"01",x"85",x"49",x"85",x"4A",x"60",x"85", -- 0x0340
    x"2F",x"60",x"A9",x"03",x"85",x"8C",x"A5",x"51", -- 0x0348
    x"F0",x"06",x"C6",x"51",x"F0",x"55",x"D0",x"52", -- 0x0350
    x"A9",x"EF",x"8D",x"20",x"91",x"AD",x"21",x"91", -- 0x0358
    x"29",x"80",x"F0",x"53",x"A9",x"DF",x"8D",x"20", -- 0x0360
    x"91",x"AD",x"21",x"91",x"29",x"01",x"D0",x"23", -- 0x0368
    x"A9",x"EF",x"8D",x"20",x"91",x"AD",x"21",x"91", -- 0x0370
    x"29",x"40",x"D0",x"17",x"A9",x"F7",x"8D",x"20", -- 0x0378
    x"91",x"AD",x"21",x"91",x"29",x"02",x"10",x"0B", -- 0x0380
    x"A2",x"77",x"BD",x"B3",x"BE",x"9D",x"78",x"14", -- 0x0388
    x"CA",x"10",x"F7",x"A9",x"FB",x"8D",x"20",x"91", -- 0x0390
    x"AD",x"21",x"91",x"29",x"80",x"D0",x"0B",x"AD", -- 0x0398
    x"00",x"90",x"18",x"69",x"01",x"29",x"0F",x"8D", -- 0x03A0
    x"00",x"90",x"60",x"A9",x"80",x"A2",x"0D",x"95", -- 0x03A8
    x"7F",x"CA",x"10",x"FB",x"4C",x"BC",x"A0",x"20", -- 0x03B0
    x"2D",x"A2",x"20",x"9F",x"A4",x"A2",x"0C",x"BD", -- 0x03B8
    x"2B",x"BF",x"9D",x"EB",x"1E",x"CA",x"10",x"F7", -- 0x03C0
    x"A9",x"16",x"85",x"51",x"A2",x"0C",x"A9",x"80", -- 0x03C8
    x"95",x"7F",x"CA",x"10",x"FB",x"60",x"A9",x"00", -- 0x03D0
    x"85",x"0B",x"A9",x"01",x"85",x"44",x"4C",x"78", -- 0x03D8
    x"AE",x"A5",x"1F",x"D0",x"7D",x"A5",x"12",x"D0", -- 0x03E0
    x"79",x"A5",x"0D",x"F0",x"1B",x"C6",x"0D",x"4A", -- 0x03E8
    x"4A",x"4A",x"8D",x"0E",x"90",x"A9",x"C8",x"8D", -- 0x03F0
    x"0A",x"90",x"A9",x"00",x"8D",x"0B",x"90",x"8D", -- 0x03F8
    x"0C",x"90",x"A9",x"80",x"8D",x"0D",x"90",x"60", -- 0x0400
    x"A5",x"0F",x"F0",x"0A",x"C6",x"0F",x"A6",x"0F", -- 0x0408
    x"BD",x"FF",x"BD",x"8D",x"0C",x"90",x"A5",x"0E", -- 0x0410
    x"F0",x"0A",x"C6",x"0E",x"A6",x"0E",x"BD",x"F3", -- 0x0418
    x"BD",x"8D",x"0C",x"90",x"A5",x"10",x"F0",x"13", -- 0x0420
    x"C6",x"10",x"D0",x"04",x"A9",x"0B",x"85",x"10", -- 0x0428
    x"A6",x"10",x"BD",x"08",x"BE",x"38",x"E5",x"13", -- 0x0430
    x"8D",x"0B",x"90",x"A9",x"00",x"8D",x"0A",x"90", -- 0x0438
    x"A5",x"11",x"F0",x"1E",x"A5",x"81",x"D0",x"1A", -- 0x0440
    x"C6",x"11",x"D0",x"16",x"E6",x"0C",x"A5",x"0C", -- 0x0448
    x"29",x"03",x"85",x"0C",x"AA",x"BD",x"EF",x"BD", -- 0x0450
    x"8D",x"0A",x"90",x"A5",x"24",x"18",x"69",x"02", -- 0x0458
    x"85",x"11",x"60",x"A9",x"00",x"85",x"0D",x"85", -- 0x0460
    x"0E",x"85",x"0F",x"85",x"10",x"85",x"12",x"8D", -- 0x0468
    x"0A",x"90",x"8D",x"0B",x"90",x"8D",x"0C",x"90", -- 0x0470
    x"8D",x"0D",x"90",x"A9",x"0F",x"8D",x"0E",x"90", -- 0x0478
    x"60",x"A9",x"00",x"85",x"0D",x"85",x"0E",x"85", -- 0x0480
    x"0F",x"85",x"10",x"8D",x"0A",x"90",x"8D",x"0B", -- 0x0488
    x"90",x"8D",x"0C",x"90",x"8D",x"0D",x"90",x"8D", -- 0x0490
    x"0E",x"90",x"A9",x"01",x"85",x"12",x"60",x"A2", -- 0x0498
    x"15",x"BD",x"EE",x"B3",x"85",x"00",x"BD",x"07", -- 0x04A0
    x"B4",x"18",x"69",x"78",x"85",x"01",x"A0",x"16", -- 0x04A8
    x"BD",x"14",x"BE",x"91",x"00",x"88",x"10",x"FB", -- 0x04B0
    x"CA",x"10",x"E6",x"A9",x"06",x"8D",x"00",x"96", -- 0x04B8
    x"8D",x"01",x"96",x"A2",x"00",x"8D",x"08",x"96", -- 0x04C0
    x"8D",x"09",x"96",x"A9",x"08",x"8D",x"0F",x"90", -- 0x04C8
    x"60",x"A9",x"02",x"A2",x"00",x"9D",x"00",x"96", -- 0x04D0
    x"9D",x"00",x"97",x"CA",x"D0",x"F7",x"60",x"A9", -- 0x04D8
    x"06",x"A2",x"00",x"9D",x"00",x"96",x"9D",x"00", -- 0x04E0
    x"97",x"CA",x"D0",x"F7",x"A9",x"19",x"8D",x"0F", -- 0x04E8
    x"90",x"60",x"8A",x"0A",x"AA",x"BD",x"13",x"B2", -- 0x04F0
    x"85",x"00",x"BD",x"14",x"B2",x"85",x"01",x"A0", -- 0x04F8
    x"00",x"B1",x"00",x"85",x"22",x"C8",x"A2",x"00", -- 0x0500
    x"B1",x"00",x"95",x"6B",x"C8",x"E8",x"E0",x"0A", -- 0x0508
    x"D0",x"F6",x"20",x"1D",x"A5",x"C6",x"22",x"F0", -- 0x0510
    x"03",x"4C",x"06",x"A5",x"60",x"98",x"48",x"A6", -- 0x0518
    x"6B",x"A5",x"6C",x"9D",x"B4",x"18",x"A9",x"00", -- 0x0520
    x"85",x"04",x"8A",x"0A",x"0A",x"26",x"04",x"0A", -- 0x0528
    x"26",x"04",x"85",x"02",x"A9",x"12",x"65",x"04", -- 0x0530
    x"85",x"03",x"A0",x"07",x"B9",x"6D",x"00",x"91", -- 0x0538
    x"02",x"88",x"10",x"F8",x"68",x"A8",x"60",x"A5", -- 0x0540
    x"24",x"D0",x"01",x"60",x"A5",x"06",x"F0",x"03", -- 0x0548
    x"4C",x"D6",x"A5",x"A5",x"19",x"30",x"04",x"A0", -- 0x0550
    x"16",x"D0",x"02",x"A0",x"00",x"A5",x"54",x"85", -- 0x0558
    x"00",x"A5",x"55",x"85",x"01",x"A9",x"05",x"85", -- 0x0560
    x"25",x"B1",x"00",x"A2",x"05",x"DD",x"21",x"B4", -- 0x0568
    x"F0",x"21",x"CA",x"10",x"F8",x"A5",x"00",x"18", -- 0x0570
    x"69",x"2E",x"90",x"02",x"E6",x"01",x"85",x"00", -- 0x0578
    x"C9",x"E3",x"A5",x"01",x"E9",x"1F",x"B0",x"04", -- 0x0580
    x"C6",x"25",x"D0",x"DD",x"A9",x"00",x"85",x"26", -- 0x0588
    x"4C",x"AB",x"A5",x"A9",x"08",x"85",x"26",x"A5", -- 0x0590
    x"19",x"49",x"FF",x"18",x"69",x"01",x"85",x"19", -- 0x0598
    x"A5",x"54",x"18",x"69",x"17",x"90",x"02",x"E6", -- 0x05A0
    x"55",x"85",x"54",x"A5",x"18",x"18",x"65",x"19", -- 0x05A8
    x"29",x"03",x"85",x"18",x"A6",x"1A",x"F0",x"06", -- 0x05B0
    x"48",x"AA",x"20",x"F2",x"A4",x"68",x"18",x"69", -- 0x05B8
    x"04",x"A6",x"1B",x"F0",x"06",x"48",x"AA",x"20", -- 0x05C0
    x"F2",x"A4",x"68",x"A6",x"1C",x"F0",x"07",x"18", -- 0x05C8
    x"69",x"04",x"AA",x"20",x"F2",x"A4",x"A5",x"06", -- 0x05D0
    x"A4",x"19",x"10",x"03",x"18",x"69",x"3C",x"A8", -- 0x05D8
    x"BE",x"27",x"B4",x"C8",x"E6",x"06",x"BD",x"78", -- 0x05E0
    x"18",x"29",x"03",x"D0",x"09",x"A5",x"06",x"C9", -- 0x05E8
    x"3C",x"D0",x"ED",x"4C",x"DB",x"A6",x"85",x"04", -- 0x05F0
    x"BD",x"3C",x"18",x"18",x"65",x"26",x"85",x"29", -- 0x05F8
    x"9D",x"3C",x"18",x"C9",x"A0",x"90",x"06",x"A9", -- 0x0600
    x"03",x"85",x"0B",x"85",x"04",x"A5",x"04",x"0A", -- 0x0608
    x"85",x"04",x"0A",x"65",x"04",x"38",x"E9",x"06", -- 0x0610
    x"85",x"27",x"BD",x"00",x"18",x"18",x"65",x"19", -- 0x0618
    x"18",x"65",x"19",x"9D",x"00",x"18",x"A5",x"18", -- 0x0620
    x"D0",x"57",x"BD",x"00",x"18",x"A4",x"19",x"30", -- 0x0628
    x"03",x"18",x"69",x"10",x"85",x"28",x"86",x"2B", -- 0x0630
    x"8A",x"18",x"65",x"19",x"AA",x"A4",x"27",x"C8", -- 0x0638
    x"BD",x"78",x"18",x"D0",x"08",x"C8",x"C8",x"C8", -- 0x0640
    x"A5",x"19",x"30",x"01",x"C8",x"98",x"20",x"E9", -- 0x0648
    x"A6",x"A6",x"2B",x"BD",x"00",x"18",x"18",x"69", -- 0x0650
    x"08",x"85",x"28",x"A5",x"27",x"20",x"E9",x"A6", -- 0x0658
    x"A5",x"27",x"18",x"69",x"04",x"85",x"04",x"BD", -- 0x0660
    x"00",x"18",x"A4",x"19",x"08",x"10",x"03",x"18", -- 0x0668
    x"69",x"10",x"85",x"28",x"A5",x"04",x"28",x"10", -- 0x0670
    x"02",x"69",x"01",x"20",x"E9",x"A6",x"4C",x"DB", -- 0x0678
    x"A6",x"A5",x"18",x"38",x"E5",x"19",x"29",x"03", -- 0x0680
    x"D0",x"34",x"8A",x"38",x"E5",x"19",x"86",x"2B", -- 0x0688
    x"AA",x"BD",x"78",x"18",x"A6",x"2B",x"29",x"03", -- 0x0690
    x"D0",x"04",x"A9",x"FA",x"D0",x"02",x"A5",x"27", -- 0x0698
    x"18",x"69",x"04",x"85",x"04",x"BD",x"00",x"18", -- 0x06A0
    x"A4",x"19",x"08",x"10",x"02",x"69",x"18",x"38", -- 0x06A8
    x"E9",x"08",x"85",x"28",x"A5",x"04",x"28",x"30", -- 0x06B0
    x"02",x"69",x"01",x"20",x"E9",x"A6",x"BD",x"00", -- 0x06B8
    x"18",x"85",x"28",x"A5",x"18",x"29",x"01",x"0A", -- 0x06C0
    x"18",x"65",x"27",x"20",x"E9",x"A6",x"A8",x"A5", -- 0x06C8
    x"28",x"18",x"69",x"08",x"85",x"28",x"C8",x"98", -- 0x06D0
    x"20",x"E9",x"A6",x"A5",x"06",x"C9",x"3C",x"D0", -- 0x06D8
    x"07",x"A9",x"00",x"85",x"06",x"4C",x"47",x"A5", -- 0x06E0
    x"60",x"48",x"84",x"2C",x"A5",x"29",x"4A",x"4A", -- 0x06E8
    x"4A",x"A8",x"B9",x"06",x"B4",x"85",x"01",x"A5", -- 0x06F0
    x"28",x"4A",x"4A",x"4A",x"18",x"79",x"ED",x"B3", -- 0x06F8
    x"90",x"02",x"E6",x"01",x"85",x"00",x"A0",x"00", -- 0x0700
    x"A9",x"20",x"91",x"00",x"68",x"48",x"C9",x"F7", -- 0x0708
    x"90",x"04",x"A9",x"20",x"D0",x"03",x"18",x"69", -- 0x0710
    x"40",x"A0",x"17",x"91",x"00",x"A4",x"2C",x"68", -- 0x0718
    x"60",x"A5",x"2F",x"48",x"29",x"07",x"18",x"69", -- 0x0720
    x"0D",x"85",x"04",x"68",x"48",x"4A",x"4A",x"4A", -- 0x0728
    x"85",x"2B",x"68",x"48",x"C5",x"08",x"F0",x"16", -- 0x0730
    x"A5",x"08",x"4A",x"4A",x"4A",x"AA",x"A9",x"20", -- 0x0738
    x"9D",x"CD",x"1F",x"9D",x"CE",x"1F",x"9D",x"CF", -- 0x0740
    x"1F",x"A6",x"04",x"20",x"F2",x"A4",x"A6",x"2B", -- 0x0748
    x"A9",x"52",x"9D",x"CD",x"1F",x"A9",x"53",x"9D", -- 0x0750
    x"CE",x"1F",x"A9",x"54",x"9D",x"CF",x"1F",x"68", -- 0x0758
    x"85",x"08",x"60",x"20",x"52",x"AC",x"A5",x"4C", -- 0x0760
    x"A6",x"2F",x"C9",x"06",x"D0",x"05",x"E0",x"98", -- 0x0768
    x"B0",x"01",x"E8",x"C9",x"04",x"D0",x"05",x"E0", -- 0x0770
    x"03",x"90",x"01",x"CA",x"86",x"2F",x"A6",x"17", -- 0x0778
    x"D0",x"11",x"A5",x"4D",x"C9",x"0A",x"D0",x"07", -- 0x0780
    x"A5",x"07",x"D0",x"07",x"4C",x"94",x"A7",x"A9", -- 0x0788
    x"00",x"85",x"07",x"60",x"A5",x"2F",x"18",x"69", -- 0x0790
    x"0E",x"85",x"5F",x"29",x"07",x"AA",x"A9",x"80", -- 0x0798
    x"CA",x"30",x"03",x"4A",x"D0",x"FA",x"A2",x"06", -- 0x07A0
    x"95",x"75",x"CA",x"10",x"FB",x"A9",x"A1",x"85", -- 0x07A8
    x"17",x"A2",x"01",x"86",x"07",x"A9",x"00",x"95", -- 0x07B0
    x"7C",x"CA",x"10",x"FB",x"85",x"63",x"85",x"6A", -- 0x07B8
    x"C6",x"3F",x"D0",x"04",x"A9",x"0F",x"85",x"3F", -- 0x07C0
    x"A9",x"09",x"85",x"0F",x"60",x"A9",x"01",x"85", -- 0x07C8
    x"80",x"A5",x"17",x"D0",x"01",x"60",x"A6",x"63", -- 0x07D0
    x"F0",x"03",x"4C",x"9A",x"A9",x"85",x"29",x"A6", -- 0x07D8
    x"5F",x"86",x"28",x"A6",x"6A",x"C9",x"A0",x"B0", -- 0x07E0
    x"0B",x"20",x"78",x"AA",x"C9",x"61",x"D0",x"04", -- 0x07E8
    x"8A",x"20",x"53",x"AA",x"A5",x"29",x"38",x"E9", -- 0x07F0
    x"08",x"C9",x"07",x"B0",x"05",x"A0",x"06",x"4C", -- 0x07F8
    x"66",x"A8",x"85",x"17",x"85",x"29",x"20",x"78", -- 0x0800
    x"AA",x"85",x"6A",x"C9",x"20",x"D0",x"19",x"E0", -- 0x0808
    x"20",x"F0",x"10",x"A9",x"21",x"85",x"6B",x"A2", -- 0x0810
    x"08",x"B5",x"75",x"95",x"6C",x"CA",x"10",x"F9", -- 0x0818
    x"20",x"1D",x"A5",x"A9",x"61",x"4C",x"53",x"AA", -- 0x0820
    x"C9",x"68",x"90",x"5F",x"C9",x"89",x"B0",x"5B", -- 0x0828
    x"38",x"E9",x"67",x"85",x"04",x"0A",x"0A",x"0A", -- 0x0830
    x"AA",x"CA",x"A5",x"29",x"A0",x"07",x"A5",x"75", -- 0x0838
    x"3D",x"40",x"13",x"D0",x"21",x"CA",x"88",x"10", -- 0x0840
    x"F5",x"A4",x"04",x"88",x"B9",x"B4",x"18",x"85", -- 0x0848
    x"04",x"E8",x"8A",x"A8",x"A2",x"00",x"B9",x"40", -- 0x0850
    x"13",x"15",x"75",x"95",x"6D",x"C8",x"E8",x"E0", -- 0x0858
    x"08",x"D0",x"F3",x"4C",x"B3",x"A8",x"84",x"04", -- 0x0860
    x"A5",x"29",x"18",x"65",x"04",x"38",x"E9",x"06", -- 0x0868
    x"85",x"29",x"85",x"17",x"A5",x"06",x"4A",x"A5", -- 0x0870
    x"28",x"E9",x"03",x"85",x"28",x"85",x"5F",x"A9", -- 0x0878
    x"00",x"A2",x"03",x"20",x"9B",x"AA",x"A9",x"06", -- 0x0880
    x"85",x"63",x"60",x"C9",x"52",x"90",x"03",x"4C", -- 0x0888
    x"63",x"A9",x"E9",x"3F",x"AA",x"BD",x"B4",x"18", -- 0x0890
    x"85",x"04",x"2D",x"D5",x"18",x"D0",x"27",x"8A", -- 0x0898
    x"0A",x"0A",x"0A",x"A8",x"A2",x"00",x"B9",x"00", -- 0x08A0
    x"12",x"15",x"75",x"95",x"6D",x"C8",x"E8",x"E0", -- 0x08A8
    x"08",x"D0",x"F3",x"A9",x"21",x"85",x"6B",x"A5", -- 0x08B0
    x"04",x"0D",x"D5",x"18",x"85",x"6C",x"20",x"1D", -- 0x08B8
    x"A5",x"A9",x"61",x"4C",x"53",x"AA",x"C6",x"29", -- 0x08C0
    x"C6",x"17",x"A5",x"28",x"4A",x"90",x"06",x"E6", -- 0x08C8
    x"28",x"A9",x"06",x"85",x"04",x"A2",x"3B",x"BD", -- 0x08D0
    x"78",x"18",x"F0",x"0E",x"BD",x"3C",x"18",x"C5", -- 0x08D8
    x"29",x"D0",x"07",x"BD",x"00",x"18",x"C5",x"28", -- 0x08E0
    x"F0",x"16",x"CA",x"10",x"EA",x"C6",x"28",x"C6", -- 0x08E8
    x"28",x"C6",x"04",x"D0",x"E0",x"A5",x"5F",x"85", -- 0x08F0
    x"28",x"E6",x"29",x"E6",x"17",x"4C",x"13",x"A8", -- 0x08F8
    x"86",x"35",x"A5",x"28",x"85",x"5F",x"4A",x"29", -- 0x0900
    x"03",x"85",x"36",x"C9",x"03",x"F0",x"14",x"69", -- 0x0908
    x"15",x"AA",x"20",x"F2",x"A4",x"A9",x"61",x"20", -- 0x0910
    x"53",x"AA",x"A0",x"01",x"A9",x"62",x"91",x"00", -- 0x0918
    x"4C",x"50",x"A9",x"86",x"2B",x"BD",x"77",x"18", -- 0x0920
    x"18",x"69",x"18",x"AA",x"20",x"F2",x"A4",x"A6", -- 0x0928
    x"2B",x"BD",x"79",x"18",x"18",x"69",x"1C",x"AA", -- 0x0930
    x"20",x"F2",x"A4",x"A2",x"20",x"20",x"F2",x"A4", -- 0x0938
    x"A9",x"61",x"20",x"53",x"AA",x"A0",x"01",x"A9", -- 0x0940
    x"62",x"91",x"00",x"C8",x"A9",x"63",x"91",x"00", -- 0x0948
    x"A6",x"35",x"BD",x"78",x"18",x"20",x"19",x"B1", -- 0x0950
    x"A9",x"86",x"85",x"63",x"85",x"81",x"A9",x"0C", -- 0x0958
    x"85",x"0E",x"60",x"C9",x"65",x"90",x"21",x"29", -- 0x0960
    x"3F",x"A8",x"B9",x"B4",x"18",x"2D",x"D5",x"18", -- 0x0968
    x"D0",x"05",x"A9",x"20",x"85",x"6B",x"60",x"A9", -- 0x0970
    x"10",x"85",x"80",x"A9",x"FF",x"85",x"43",x"A9", -- 0x0978
    x"00",x"85",x"17",x"A9",x"18",x"85",x"13",x"60", -- 0x0980
    x"38",x"E9",x"55",x"4A",x"4A",x"AA",x"B5",x"60", -- 0x0988
    x"C9",x"05",x"90",x"01",x"60",x"A0",x"00",x"4C", -- 0x0990
    x"66",x"A8",x"A5",x"5F",x"85",x"28",x"A5",x"17", -- 0x0998
    x"85",x"29",x"C6",x"63",x"30",x"0D",x"F0",x"01", -- 0x09A0
    x"60",x"A2",x"03",x"20",x"E9",x"AB",x"A9",x"00", -- 0x09A8
    x"85",x"17",x"60",x"A5",x"63",x"C9",x"81",x"F0", -- 0x09B0
    x"03",x"4C",x"52",x"AA",x"A0",x"00",x"A5",x"36", -- 0x09B8
    x"C9",x"03",x"F0",x"08",x"A9",x"20",x"20",x"53", -- 0x09C0
    x"AA",x"4C",x"16",x"AA",x"A5",x"06",x"A4",x"19", -- 0x09C8
    x"10",x"03",x"18",x"69",x"3C",x"A8",x"BE",x"27", -- 0x09D0
    x"B4",x"E4",x"35",x"D0",x"0B",x"A9",x"20",x"20", -- 0x09D8
    x"53",x"AA",x"A0",x"01",x"91",x"00",x"D0",x"2E", -- 0x09E0
    x"A0",x"00",x"A6",x"35",x"BD",x"77",x"18",x"D0", -- 0x09E8
    x"04",x"A9",x"20",x"D0",x"08",x"0A",x"85",x"04", -- 0x09F0
    x"0A",x"65",x"04",x"69",x"3F",x"20",x"53",x"AA", -- 0x09F8
    x"C8",x"A9",x"20",x"91",x"00",x"BD",x"79",x"18", -- 0x0A00
    x"D0",x"04",x"A9",x"20",x"D0",x"08",x"0A",x"85", -- 0x0A08
    x"04",x"0A",x"65",x"04",x"69",x"3E",x"C8",x"91", -- 0x0A10
    x"00",x"A6",x"35",x"A9",x"00",x"9D",x"78",x"18", -- 0x0A18
    x"A5",x"87",x"29",x"80",x"49",x"80",x"85",x"81", -- 0x0A20
    x"C6",x"24",x"A5",x"24",x"C9",x"08",x"90",x"03", -- 0x0A28
    x"4C",x"AE",x"A9",x"A2",x"00",x"86",x"1A",x"86", -- 0x0A30
    x"1B",x"86",x"1C",x"E8",x"86",x"4B",x"A0",x"3B", -- 0x0A38
    x"B9",x"78",x"18",x"F0",x"03",x"AA",x"95",x"19", -- 0x0A40
    x"88",x"10",x"F5",x"A9",x"80",x"85",x"86",x"4C", -- 0x0A48
    x"AE",x"A9",x"60",x"84",x"2C",x"48",x"A5",x"29", -- 0x0A50
    x"4A",x"4A",x"4A",x"A8",x"B9",x"07",x"B4",x"85", -- 0x0A58
    x"01",x"A5",x"28",x"4A",x"4A",x"4A",x"18",x"79", -- 0x0A60
    x"EE",x"B3",x"90",x"02",x"E6",x"01",x"85",x"00", -- 0x0A68
    x"A0",x"00",x"68",x"91",x"00",x"A4",x"2C",x"60", -- 0x0A70
    x"84",x"2C",x"A5",x"29",x"4A",x"4A",x"4A",x"A8", -- 0x0A78
    x"B9",x"07",x"B4",x"85",x"01",x"A5",x"28",x"4A", -- 0x0A80
    x"4A",x"4A",x"18",x"79",x"EE",x"B3",x"90",x"02", -- 0x0A88
    x"E6",x"01",x"85",x"00",x"A0",x"00",x"B1",x"00", -- 0x0A90
    x"A4",x"2C",x"60",x"8A",x"85",x"30",x"0A",x"0A", -- 0x0A98
    x"AA",x"85",x"31",x"20",x"78",x"AA",x"95",x"8E", -- 0x0AA0
    x"A0",x"17",x"B1",x"00",x"95",x"8F",x"A0",x"01", -- 0x0AA8
    x"B1",x"00",x"95",x"90",x"A0",x"18",x"B1",x"00", -- 0x0AB0
    x"95",x"91",x"A2",x"1F",x"A9",x"00",x"95",x"9E", -- 0x0AB8
    x"CA",x"10",x"FB",x"A5",x"28",x"29",x"07",x"0A", -- 0x0AC0
    x"0A",x"0A",x"A6",x"30",x"E0",x"03",x"F0",x"04", -- 0x0AC8
    x"09",x"80",x"D0",x"01",x"0A",x"A8",x"A5",x"29", -- 0x0AD0
    x"29",x"07",x"AA",x"A9",x"08",x"85",x"04",x"B9", -- 0x0AD8
    x"E4",x"B5",x"95",x"9E",x"B9",x"EC",x"B5",x"95", -- 0x0AE0
    x"AE",x"E8",x"C8",x"C6",x"04",x"D0",x"F0",x"A9", -- 0x0AE8
    x"03",x"85",x"32",x"A5",x"32",x"05",x"31",x"AA", -- 0x0AF0
    x"A9",x"04",x"85",x"50",x"B5",x"8E",x"C9",x"68", -- 0x0AF8
    x"90",x"68",x"C9",x"89",x"B0",x"64",x"38",x"E9", -- 0x0B00
    x"40",x"85",x"34",x"8A",x"18",x"69",x"15",x"85", -- 0x0B08
    x"6B",x"85",x"4F",x"A5",x"34",x"38",x"E9",x"28", -- 0x0B10
    x"0A",x"0A",x"0A",x"AA",x"86",x"2B",x"A5",x"32", -- 0x0B18
    x"0A",x"0A",x"0A",x"A8",x"84",x"2C",x"A9",x"08", -- 0x0B20
    x"85",x"04",x"B9",x"9E",x"00",x"1D",x"40",x"13", -- 0x0B28
    x"48",x"E8",x"C8",x"C6",x"04",x"D0",x"F3",x"A2", -- 0x0B30
    x"07",x"68",x"95",x"6D",x"CA",x"10",x"FA",x"20", -- 0x0B38
    x"1D",x"A5",x"A6",x"2B",x"A4",x"2C",x"A9",x"08", -- 0x0B40
    x"85",x"04",x"B9",x"9E",x"00",x"49",x"FF",x"3D", -- 0x0B48
    x"40",x"13",x"9D",x"40",x"13",x"48",x"E8",x"C8", -- 0x0B50
    x"C6",x"04",x"D0",x"EE",x"A2",x"07",x"68",x"95", -- 0x0B58
    x"6D",x"CA",x"10",x"FA",x"A5",x"34",x"85",x"6B", -- 0x0B60
    x"D0",x"68",x"C9",x"55",x"90",x"46",x"C9",x"65", -- 0x0B68
    x"B0",x"42",x"48",x"38",x"E5",x"31",x"C9",x"55", -- 0x0B70
    x"F0",x"36",x"C9",x"56",x"F0",x"32",x"C9",x"57", -- 0x0B78
    x"F0",x"2E",x"C9",x"58",x"F0",x"2A",x"68",x"38", -- 0x0B80
    x"E9",x"55",x"A8",x"4A",x"4A",x"AA",x"B5",x"60", -- 0x0B88
    x"F0",x"22",x"A5",x"32",x"05",x"31",x"AA",x"B9", -- 0x0B90
    x"8E",x"00",x"95",x"8E",x"84",x"04",x"A6",x"04", -- 0x0B98
    x"C6",x"50",x"D0",x"09",x"A5",x"32",x"05",x"31", -- 0x0BA0
    x"AA",x"A9",x"20",x"95",x"8E",x"4C",x"FE",x"AA", -- 0x0BA8
    x"68",x"4C",x"A4",x"AB",x"A5",x"32",x"48",x"0A", -- 0x0BB0
    x"0A",x"0A",x"AA",x"A0",x"00",x"B5",x"9E",x"99", -- 0x0BB8
    x"6D",x"00",x"E8",x"C8",x"C0",x"08",x"D0",x"F5", -- 0x0BC0
    x"68",x"05",x"31",x"18",x"69",x"15",x"85",x"6B", -- 0x0BC8
    x"85",x"4F",x"20",x"1D",x"A5",x"A6",x"32",x"BC", -- 0x0BD0
    x"44",x"B7",x"A5",x"4F",x"18",x"69",x"40",x"91", -- 0x0BD8
    x"00",x"C6",x"32",x"30",x"03",x"4C",x"F3",x"AA", -- 0x0BE0
    x"60",x"8A",x"0A",x"0A",x"AA",x"18",x"69",x"55", -- 0x0BE8
    x"85",x"04",x"A0",x"00",x"20",x"78",x"AA",x"C5", -- 0x0BF0
    x"04",x"D0",x"0E",x"B5",x"8E",x"C9",x"52",x"90", -- 0x0BF8
    x"06",x"C9",x"65",x"B0",x"02",x"A9",x"20",x"91", -- 0x0C00
    x"00",x"A0",x"17",x"E6",x"04",x"B1",x"00",x"C5", -- 0x0C08
    x"04",x"D0",x"0E",x"B5",x"8F",x"C9",x"52",x"90", -- 0x0C10
    x"06",x"C9",x"65",x"B0",x"02",x"A9",x"20",x"91", -- 0x0C18
    x"00",x"A0",x"01",x"E6",x"04",x"B1",x"00",x"C5", -- 0x0C20
    x"04",x"D0",x"0E",x"B5",x"90",x"C9",x"52",x"90", -- 0x0C28
    x"06",x"C9",x"65",x"B0",x"02",x"A9",x"20",x"91", -- 0x0C30
    x"00",x"A0",x"18",x"E6",x"04",x"B1",x"00",x"C5", -- 0x0C38
    x"04",x"D0",x"0E",x"B5",x"91",x"C9",x"52",x"90", -- 0x0C40
    x"06",x"C9",x"65",x"B0",x"02",x"A9",x"20",x"91", -- 0x0C48
    x"00",x"60",x"A9",x"00",x"85",x"4D",x"85",x"4C", -- 0x0C50
    x"A2",x"03",x"BD",x"CB",x"AC",x"8D",x"20",x"91", -- 0x0C58
    x"AD",x"21",x"91",x"CD",x"21",x"91",x"D0",x"F8", -- 0x0C60
    x"3D",x"CF",x"AC",x"D0",x"05",x"BD",x"D3",x"AC", -- 0x0C68
    x"85",x"4C",x"CA",x"10",x"E5",x"A2",x"01",x"A9", -- 0x0C70
    x"FB",x"8D",x"20",x"91",x"AD",x"21",x"91",x"CD", -- 0x0C78
    x"21",x"91",x"D0",x"F8",x"3D",x"D7",x"AC",x"D0", -- 0x0C80
    x"05",x"BD",x"D9",x"AC",x"85",x"4D",x"CA",x"10", -- 0x0C88
    x"E6",x"A2",x"7F",x"8E",x"22",x"91",x"AD",x"20", -- 0x0C90
    x"91",x"CD",x"20",x"91",x"D0",x"F8",x"A2",x"FF", -- 0x0C98
    x"8E",x"22",x"91",x"A2",x"7F",x"8E",x"20",x"91", -- 0x0CA0
    x"29",x"80",x"D0",x"04",x"A9",x"06",x"85",x"4C", -- 0x0CA8
    x"AD",x"1F",x"91",x"CD",x"1F",x"91",x"D0",x"F8", -- 0x0CB0
    x"A8",x"29",x"10",x"D0",x"04",x"A9",x"04",x"85", -- 0x0CB8
    x"4C",x"98",x"29",x"20",x"D0",x"04",x"A9",x"0A", -- 0x0CC0
    x"85",x"4D",x"60",x"EF",x"FB",x"FB",x"FD",x"20", -- 0x0CC8
    x"20",x"40",x"20",x"02",x"04",x"06",x"08",x"02", -- 0x0CD0
    x"04",x"0A",x"0D",x"A9",x"03",x"85",x"85",x"A6", -- 0x0CD8
    x"4B",x"B5",x"14",x"F0",x"04",x"CA",x"10",x"F9", -- 0x0CE0
    x"60",x"86",x"2B",x"A4",x"09",x"BE",x"11",x"BA", -- 0x0CE8
    x"18",x"BD",x"78",x"18",x"D0",x"0B",x"8A",x"69", -- 0x0CF0
    x"0C",x"AA",x"C9",x"3C",x"E6",x"09",x"90",x"F1", -- 0x0CF8
    x"60",x"8A",x"A8",x"A6",x"2B",x"B9",x"00",x"18", -- 0x0D00
    x"29",x"06",x"C9",x"02",x"D0",x"01",x"60",x"4A", -- 0x0D08
    x"84",x"2C",x"A8",x"B9",x"48",x"B7",x"95",x"56", -- 0x0D10
    x"A4",x"2C",x"B9",x"3C",x"18",x"18",x"69",x"0C", -- 0x0D18
    x"95",x"14",x"85",x"29",x"A9",x"00",x"95",x"60", -- 0x0D20
    x"B9",x"00",x"18",x"18",x"69",x"04",x"95",x"5C", -- 0x0D28
    x"85",x"28",x"A0",x"17",x"20",x"1B",x"B0",x"B1", -- 0x0D30
    x"00",x"C9",x"55",x"90",x"09",x"C9",x"61",x"B0", -- 0x0D38
    x"05",x"A9",x"00",x"95",x"14",x"60",x"A5",x"28", -- 0x0D40
    x"29",x"06",x"0A",x"0A",x"0A",x"0A",x"0A",x"85", -- 0x0D48
    x"04",x"BD",x"0B",x"BA",x"18",x"65",x"04",x"85", -- 0x0D50
    x"00",x"BD",x"0E",x"BA",x"69",x"00",x"85",x"01", -- 0x0D58
    x"E8",x"A0",x"3F",x"8A",x"0A",x"06",x"2B",x"0A", -- 0x0D60
    x"0A",x"0A",x"0A",x"0A",x"AA",x"CA",x"B1",x"00", -- 0x0D68
    x"9D",x"34",x"19",x"CA",x"88",x"10",x"F7",x"A6", -- 0x0D70
    x"2B",x"20",x"78",x"AA",x"95",x"64",x"A0",x"17", -- 0x0D78
    x"B1",x"00",x"95",x"65",x"60",x"A9",x"02",x"85", -- 0x0D80
    x"38",x"A9",x"03",x"85",x"7F",x"A5",x"38",x"AA", -- 0x0D88
    x"0A",x"85",x"39",x"0A",x"85",x"3A",x"0A",x"0A", -- 0x0D90
    x"0A",x"0A",x"85",x"3B",x"B5",x"5C",x"85",x"28", -- 0x0D98
    x"B5",x"14",x"85",x"29",x"D0",x"03",x"4C",x"01", -- 0x0DA0
    x"B0",x"B5",x"60",x"F0",x"03",x"4C",x"09",x"B0", -- 0x0DA8
    x"A5",x"3A",x"18",x"69",x"55",x"85",x"04",x"A6", -- 0x0DB0
    x"39",x"A0",x"00",x"20",x"78",x"AA",x"C5",x"04", -- 0x0DB8
    x"D0",x"0E",x"B5",x"64",x"C9",x"55",x"90",x"06", -- 0x0DC0
    x"C9",x"65",x"B0",x"02",x"90",x"02",x"91",x"00", -- 0x0DC8
    x"E6",x"04",x"A0",x"17",x"B1",x"00",x"C5",x"04", -- 0x0DD0
    x"D0",x"0E",x"B5",x"65",x"C9",x"55",x"90",x"06", -- 0x0DD8
    x"C9",x"65",x"B0",x"02",x"90",x"02",x"91",x"00", -- 0x0DE0
    x"A5",x"29",x"18",x"69",x"04",x"85",x"29",x"A6", -- 0x0DE8
    x"38",x"95",x"14",x"C9",x"A8",x"90",x"03",x"4C", -- 0x0DF0
    x"85",x"AF",x"A9",x"00",x"85",x"3C",x"85",x"3D", -- 0x0DF8
    x"85",x"3E",x"20",x"1B",x"B0",x"A4",x"3E",x"A5", -- 0x0E00
    x"3C",x"05",x"39",x"AA",x"B1",x"00",x"95",x"64", -- 0x0E08
    x"C9",x"20",x"D0",x"3B",x"A5",x"29",x"29",x"0C", -- 0x0E10
    x"0A",x"0A",x"05",x"3B",x"05",x"3D",x"A8",x"A5", -- 0x0E18
    x"3A",x"18",x"69",x"15",x"65",x"3C",x"85",x"6B", -- 0x0E20
    x"18",x"69",x"40",x"85",x"33",x"A6",x"38",x"B5", -- 0x0E28
    x"56",x"85",x"6C",x"A2",x"00",x"B9",x"34",x"19", -- 0x0E30
    x"95",x"6D",x"C8",x"E8",x"E0",x"08",x"D0",x"F5", -- 0x0E38
    x"20",x"1D",x"A5",x"20",x"1B",x"B0",x"A5",x"33", -- 0x0E40
    x"A4",x"3E",x"91",x"00",x"4C",x"E8",x"AF",x"C9", -- 0x0E48
    x"55",x"90",x"03",x"4C",x"EE",x"AE",x"38",x"E9", -- 0x0E50
    x"40",x"A8",x"A6",x"38",x"B9",x"B4",x"18",x"35", -- 0x0E58
    x"56",x"F0",x"42",x"C0",x"12",x"90",x"3B",x"84", -- 0x0E60
    x"0A",x"A9",x"20",x"20",x"53",x"AA",x"A0",x"17", -- 0x0E68
    x"91",x"00",x"A6",x"38",x"A9",x"00",x"95",x"14", -- 0x0E70
    x"A9",x"80",x"A2",x"05",x"95",x"81",x"CA",x"10", -- 0x0E78
    x"FB",x"85",x"8B",x"A9",x"00",x"85",x"87",x"85", -- 0x0E80
    x"0A",x"A5",x"2F",x"4A",x"29",x"03",x"85",x"46", -- 0x0E88
    x"A9",x"0F",x"85",x"45",x"A9",x"7F",x"85",x"0D", -- 0x0E90
    x"A5",x"1F",x"D0",x"03",x"20",x"D1",x"A4",x"4C", -- 0x0E98
    x"01",x"B0",x"4C",x"85",x"AF",x"84",x"04",x"A6", -- 0x0EA0
    x"38",x"B9",x"B4",x"18",x"15",x"56",x"85",x"6C", -- 0x0EA8
    x"A5",x"29",x"29",x"0C",x"0A",x"0A",x"05",x"3B", -- 0x0EB0
    x"05",x"3D",x"A8",x"A5",x"3A",x"18",x"69",x"15", -- 0x0EB8
    x"65",x"3C",x"85",x"6B",x"18",x"69",x"40",x"85", -- 0x0EC0
    x"33",x"A5",x"04",x"0A",x"0A",x"0A",x"AA",x"A9", -- 0x0EC8
    x"08",x"85",x"34",x"B9",x"34",x"19",x"1D",x"00", -- 0x0ED0
    x"12",x"48",x"E8",x"C8",x"C6",x"34",x"D0",x"F3", -- 0x0ED8
    x"A2",x"07",x"68",x"95",x"6D",x"CA",x"10",x"FA", -- 0x0EE0
    x"4C",x"40",x"AE",x"4C",x"A3",x"AF",x"C9",x"68", -- 0x0EE8
    x"90",x"F9",x"C9",x"89",x"B0",x"F5",x"38",x"E9", -- 0x0EF0
    x"68",x"0A",x"0A",x"0A",x"A8",x"A6",x"38",x"A9", -- 0x0EF8
    x"07",x"85",x"04",x"B9",x"40",x"13",x"35",x"56", -- 0x0F00
    x"D0",x"3E",x"C8",x"C6",x"04",x"10",x"F4",x"A5", -- 0x0F08
    x"29",x"29",x"0C",x"0A",x"0A",x"05",x"3B",x"05", -- 0x0F10
    x"3D",x"AA",x"A5",x"3A",x"18",x"69",x"15",x"65", -- 0x0F18
    x"3C",x"85",x"6B",x"18",x"69",x"40",x"85",x"33", -- 0x0F20
    x"98",x"E9",x"07",x"A8",x"A9",x"08",x"85",x"34", -- 0x0F28
    x"BD",x"34",x"19",x"19",x"40",x"13",x"48",x"E8", -- 0x0F30
    x"C8",x"C6",x"34",x"D0",x"F3",x"A2",x"07",x"68", -- 0x0F38
    x"95",x"6D",x"CA",x"10",x"FA",x"4C",x"40",x"AE", -- 0x0F40
    x"A5",x"3E",x"F0",x"15",x"20",x"1B",x"B0",x"A6", -- 0x0F48
    x"39",x"A0",x"00",x"B5",x"64",x"C9",x"52",x"90", -- 0x0F50
    x"06",x"C9",x"65",x"B0",x"02",x"A9",x"20",x"91", -- 0x0F58
    x"00",x"A6",x"38",x"A5",x"29",x"18",x"69",x"02", -- 0x0F60
    x"65",x"3D",x"E5",x"04",x"85",x"29",x"95",x"14", -- 0x0F68
    x"A5",x"28",x"38",x"E9",x"04",x"85",x"28",x"95", -- 0x0F70
    x"5C",x"A9",x"06",x"95",x"60",x"A6",x"38",x"20", -- 0x0F78
    x"9B",x"AA",x"4C",x"01",x"B0",x"A5",x"3E",x"F0", -- 0x0F80
    x"15",x"20",x"1B",x"B0",x"A6",x"39",x"B5",x"64", -- 0x0F88
    x"C9",x"52",x"90",x"06",x"C9",x"65",x"B0",x"02", -- 0x0F90
    x"A9",x"20",x"A0",x"00",x"91",x"00",x"A6",x"38", -- 0x0F98
    x"4C",x"70",x"AF",x"C9",x"61",x"B0",x"28",x"38", -- 0x0FA0
    x"E9",x"55",x"4A",x"4A",x"AA",x"B5",x"60",x"F0", -- 0x0FA8
    x"12",x"A4",x"3E",x"F0",x"05",x"A9",x"20",x"20", -- 0x0FB0
    x"53",x"AA",x"A6",x"38",x"A9",x"00",x"95",x"14", -- 0x0FB8
    x"4C",x"01",x"B0",x"A5",x"3C",x"05",x"39",x"AA", -- 0x0FC0
    x"A9",x"20",x"95",x"64",x"4C",x"14",x"AE",x"C9", -- 0x0FC8
    x"65",x"B0",x"12",x"A5",x"63",x"D0",x"03",x"4C", -- 0x0FD0
    x"85",x"AF",x"A5",x"09",x"4A",x"4A",x"90",x"08", -- 0x0FD8
    x"4A",x"90",x"05",x"B0",x"A0",x"4C",x"85",x"AF", -- 0x0FE0
    x"A5",x"3C",x"D0",x"15",x"A5",x"29",x"29",x"07", -- 0x0FE8
    x"F0",x"0F",x"A9",x"01",x"85",x"3C",x"A9",x"08", -- 0x0FF0
    x"85",x"3D",x"A9",x"17",x"85",x"3E",x"4C",x"02", -- 0x0FF8
    x"AE",x"C6",x"38",x"30",x"03",x"4C",x"8D",x"AD", -- 0x1000
    x"60",x"D6",x"60",x"D0",x"0B",x"A6",x"38",x"20", -- 0x1008
    x"E9",x"AB",x"A6",x"38",x"A9",x"00",x"95",x"14", -- 0x1010
    x"4C",x"01",x"B0",x"84",x"2C",x"A5",x"29",x"4A", -- 0x1018
    x"4A",x"4A",x"A8",x"B9",x"07",x"B4",x"85",x"01", -- 0x1020
    x"A5",x"28",x"4A",x"4A",x"4A",x"18",x"79",x"EE", -- 0x1028
    x"B3",x"90",x"02",x"E6",x"01",x"85",x"00",x"A4", -- 0x1030
    x"2C",x"60",x"A9",x"7F",x"85",x"86",x"C6",x"40", -- 0x1038
    x"30",x"01",x"60",x"A9",x"0B",x"85",x"40",x"A5", -- 0x1040
    x"3F",x"4A",x"4A",x"90",x"08",x"A9",x"00",x"85", -- 0x1048
    x"41",x"A9",x"02",x"D0",x"06",x"A9",x"A8",x"85", -- 0x1050
    x"41",x"A9",x"FE",x"85",x"42",x"A9",x"00",x"85", -- 0x1058
    x"43",x"85",x"83",x"A9",x"0C",x"85",x"10",x"60", -- 0x1060
    x"A9",x"03",x"85",x"83",x"A5",x"43",x"10",x"4C", -- 0x1068
    x"C9",x"FF",x"D0",x"0F",x"A9",x"87",x"85",x"43", -- 0x1070
    x"A5",x"41",x"4A",x"29",x"03",x"69",x"26",x"AA", -- 0x1078
    x"4C",x"F2",x"A4",x"C6",x"43",x"10",x"01",x"60", -- 0x1080
    x"A5",x"41",x"4A",x"4A",x"4A",x"A8",x"A6",x"3F", -- 0x1088
    x"BD",x"08",x"BC",x"48",x"4A",x"4A",x"4A",x"4A", -- 0x1090
    x"F0",x"06",x"09",x"30",x"99",x"17",x"1E",x"C8", -- 0x1098
    x"68",x"48",x"29",x"0F",x"09",x"30",x"99",x"17", -- 0x10A0
    x"1E",x"A9",x"30",x"99",x"18",x"1E",x"A9",x"20", -- 0x10A8
    x"99",x"19",x"1E",x"68",x"20",x"19",x"B1",x"A9", -- 0x10B0
    x"14",x"85",x"43",x"60",x"F0",x"11",x"C6",x"43", -- 0x10B8
    x"F0",x"01",x"60",x"A5",x"41",x"A2",x"FC",x"86", -- 0x10C0
    x"41",x"A2",x"00",x"86",x"13",x"F0",x"02",x"A5", -- 0x10C8
    x"41",x"4A",x"4A",x"4A",x"A8",x"A9",x"20",x"99", -- 0x10D0
    x"17",x"1E",x"99",x"18",x"1E",x"99",x"19",x"1E", -- 0x10D8
    x"A5",x"41",x"18",x"65",x"42",x"85",x"41",x"C9", -- 0x10E0
    x"AA",x"90",x"0C",x"A9",x"80",x"85",x"83",x"A9", -- 0x10E8
    x"00",x"85",x"10",x"8D",x"0B",x"90",x"60",x"4A", -- 0x10F0
    x"48",x"4A",x"4A",x"85",x"2C",x"68",x"29",x"03", -- 0x10F8
    x"18",x"69",x"22",x"AA",x"20",x"F2",x"A4",x"A4", -- 0x1100
    x"2C",x"A9",x"65",x"99",x"17",x"1E",x"A9",x"66", -- 0x1108
    x"99",x"18",x"1E",x"A9",x"67",x"99",x"19",x"1E", -- 0x1110
    x"60",x"F8",x"18",x"65",x"20",x"85",x"20",x"A5", -- 0x1118
    x"21",x"69",x"00",x"85",x"21",x"D8",x"F0",x"11", -- 0x1120
    x"A5",x"20",x"C9",x"50",x"90",x"0B",x"A6",x"1E", -- 0x1128
    x"D0",x"07",x"E6",x"44",x"20",x"EA",x"B1",x"85", -- 0x1130
    x"1E",x"A9",x"30",x"8D",x"06",x"1E",x"A9",x"20", -- 0x1138
    x"8D",x"07",x"1E",x"A5",x"1F",x"D0",x"1A",x"A2", -- 0x1140
    x"00",x"A5",x"21",x"20",x"50",x"B1",x"A5",x"20", -- 0x1148
    x"48",x"4A",x"4A",x"4A",x"4A",x"20",x"5B",x"B1", -- 0x1150
    x"68",x"29",x"0F",x"09",x"30",x"9D",x"02",x"1E", -- 0x1158
    x"E8",x"60",x"A9",x"06",x"85",x"87",x"A5",x"2F", -- 0x1160
    x"4A",x"4A",x"4A",x"AA",x"C6",x"45",x"30",x"24", -- 0x1168
    x"A9",x"20",x"9D",x"CC",x"1F",x"9D",x"D0",x"1F", -- 0x1170
    x"A9",x"52",x"9D",x"CD",x"1F",x"A9",x"53",x"9D", -- 0x1178
    x"CE",x"1F",x"A9",x"54",x"9D",x"CF",x"1F",x"A5", -- 0x1180
    x"46",x"49",x"04",x"85",x"46",x"18",x"69",x"2A", -- 0x1188
    x"AA",x"4C",x"F2",x"A4",x"A9",x"20",x"9D",x"CD", -- 0x1190
    x"1F",x"9D",x"CE",x"1F",x"9D",x"CF",x"1F",x"A5", -- 0x1198
    x"1F",x"F0",x"02",x"85",x"44",x"C6",x"44",x"20", -- 0x11A0
    x"EA",x"B1",x"A2",x"09",x"BD",x"3A",x"B7",x"95", -- 0x11A8
    x"7F",x"CA",x"10",x"F8",x"A5",x"41",x"C9",x"A9", -- 0x11B0
    x"90",x"04",x"A9",x"80",x"85",x"83",x"A2",x"03", -- 0x11B8
    x"86",x"2F",x"CA",x"86",x"08",x"A9",x"00",x"85", -- 0x11C0
    x"0D",x"85",x"0E",x"85",x"0F",x"8D",x"0A",x"90", -- 0x11C8
    x"8D",x"0D",x"90",x"A9",x"0F",x"8D",x"0E",x"90", -- 0x11D0
    x"20",x"9F",x"A4",x"A5",x"24",x"C9",x"08",x"B0", -- 0x11D8
    x"04",x"A9",x"80",x"85",x"86",x"A2",x"32",x"4C", -- 0x11E0
    x"F2",x"A4",x"A2",x"05",x"A9",x"20",x"9D",x"11", -- 0x11E8
    x"1E",x"CA",x"10",x"FA",x"A5",x"44",x"48",x"09", -- 0x11F0
    x"30",x"8D",x"10",x"1E",x"68",x"0A",x"AA",x"D0", -- 0x11F8
    x"01",x"60",x"CA",x"CA",x"D0",x"01",x"60",x"A9", -- 0x1200
    x"8B",x"9D",x"10",x"1E",x"A9",x"8A",x"9D",x"0F", -- 0x1208
    x"1E",x"D0",x"EF",x"79",x"B2",x"B8",x"B2",x"A3", -- 0x1210
    x"B2",x"8E",x"B2",x"CD",x"B2",x"E2",x"B2",x"F7", -- 0x1218
    x"B2",x"0C",x"B3",x"21",x"B3",x"36",x"B3",x"4B", -- 0x1220
    x"B3",x"60",x"B3",x"75",x"B3",x"00",x"B5",x"1F", -- 0x1228
    x"B5",x"34",x"B5",x"49",x"B5",x"68",x"B5",x"87", -- 0x1230
    x"B5",x"A6",x"B5",x"C5",x"B5",x"A4",x"B6",x"B9", -- 0x1238
    x"B6",x"CE",x"B6",x"E3",x"B6",x"EE",x"B6",x"F9", -- 0x1240
    x"B6",x"E3",x"B6",x"04",x"B7",x"0F",x"B7",x"1A", -- 0x1248
    x"B7",x"04",x"B7",x"25",x"B7",x"6B",x"B7",x"11", -- 0x1250
    x"BB",x"30",x"BB",x"4F",x"BB",x"6E",x"BB",x"8D", -- 0x1258
    x"BB",x"AC",x"BB",x"CB",x"BB",x"EA",x"BB",x"18", -- 0x1260
    x"BC",x"37",x"BC",x"56",x"BC",x"75",x"BC",x"94", -- 0x1268
    x"BC",x"B3",x"BC",x"D2",x"BC",x"F1",x"BC",x"10", -- 0x1270
    x"BD",x"02",x"00",x"FF",x"3C",x"FF",x"FF",x"99", -- 0x1278
    x"FF",x"E7",x"99",x"C3",x"01",x"C3",x"00",x"81", -- 0x1280
    x"C3",x"C3",x"C3",x"00",x"81",x"00",x"02",x"02", -- 0x1288
    x"0F",x"00",x"07",x"0F",x"0E",x"0F",x"01",x"03", -- 0x1290
    x"0C",x"03",x"FF",x"F0",x"FE",x"FF",x"67",x"FF", -- 0x1298
    x"98",x"6C",x"03",x"02",x"00",x"3F",x"03",x"1F", -- 0x12A0
    x"3F",x"39",x"3F",x"0E",x"19",x"0C",x"01",x"FC", -- 0x12A8
    x"C0",x"F8",x"FC",x"9C",x"FC",x"70",x"98",x"30", -- 0x12B0
    x"02",x"02",x"FF",x"0F",x"7F",x"FF",x"E6",x"FF", -- 0x12B8
    x"19",x"36",x"C0",x"03",x"F0",x"00",x"E0",x"F0", -- 0x12C0
    x"70",x"F0",x"80",x"C0",x"30",x"02",x"06",x"FF", -- 0x12C8
    x"41",x"22",x"7F",x"DD",x"FF",x"7F",x"41",x"36", -- 0x12D0
    x"07",x"C1",x"00",x"00",x"00",x"80",x"C1",x"41", -- 0x12D8
    x"41",x"00",x"02",x"08",x"FF",x"10",x"48",x"5F", -- 0x12E0
    x"77",x"3F",x"1F",x"10",x"20",x"09",x"F0",x"40", -- 0x12E8
    x"90",x"D0",x"70",x"E0",x"C0",x"40",x"20",x"02", -- 0x12F0
    x"06",x"1F",x"04",x"02",x"07",x"0D",x"1F",x"17", -- 0x12F8
    x"14",x"03",x"07",x"FC",x"10",x"20",x"F0",x"D8", -- 0x1300
    x"FC",x"F4",x"14",x"60",x"02",x"08",x"07",x"01", -- 0x1308
    x"04",x"05",x"07",x"03",x"01",x"01",x"02",x"09", -- 0x1310
    x"FF",x"04",x"89",x"FD",x"77",x"FE",x"FC",x"04", -- 0x1318
    x"02",x"02",x"0C",x"FF",x"18",x"3C",x"7E",x"DB", -- 0x1320
    x"FF",x"5A",x"81",x"42",x"0D",x"00",x"00",x"00", -- 0x1328
    x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"0E", -- 0x1330
    x"3F",x"06",x"0F",x"1F",x"36",x"3F",x"09",x"16", -- 0x1338
    x"29",x"0F",x"C0",x"00",x"00",x"80",x"C0",x"C0", -- 0x1340
    x"00",x"80",x"40",x"02",x"0C",x"0F",x"01",x"03", -- 0x1348
    x"07",x"0D",x"0F",x"05",x"08",x"04",x"0D",x"F0", -- 0x1350
    x"80",x"C0",x"E0",x"B0",x"F0",x"A0",x"10",x"20", -- 0x1358
    x"02",x"0E",x"03",x"00",x"00",x"01",x"03",x"03", -- 0x1360
    x"00",x"01",x"02",x"0F",x"FC",x"60",x"F0",x"F8", -- 0x1368
    x"6C",x"FC",x"90",x"68",x"94",x"0C",x"04",x"03", -- 0x1370
    x"00",x"01",x"03",x"03",x"03",x"00",x"01",x"00", -- 0x1378
    x"05",x"C0",x"00",x"80",x"C0",x"C0",x"C0",x"00", -- 0x1380
    x"80",x"00",x"0A",x"01",x"00",x"00",x"00",x"00", -- 0x1388
    x"01",x"01",x"01",x"00",x"0B",x"C0",x"00",x"00", -- 0x1390
    x"00",x"80",x"C0",x"40",x"40",x"00",x"10",x"00", -- 0x1398
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13A0
    x"11",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13A8
    x"00",x"00",x"14",x"00",x"00",x"00",x"00",x"00", -- 0x13B0
    x"00",x"00",x"00",x"00",x"4A",x"FF",x"02",x"07", -- 0x13B8
    x"07",x"7F",x"FF",x"FF",x"FF",x"FF",x"4B",x"F8", -- 0x13C0
    x"00",x"00",x"00",x"F0",x"F8",x"F8",x"F8",x"F8", -- 0x13C8
    x"4C",x"01",x"BF",x"BF",x"BF",x"BF",x"BF",x"BF", -- 0x13D0
    x"81",x"FF",x"4D",x"01",x"E7",x"DB",x"BD",x"81", -- 0x13D8
    x"BD",x"BD",x"BD",x"FF",x"4E",x"01",x"FF",x"FF", -- 0x13E0
    x"F7",x"FF",x"FF",x"F7",x"F7",x"EF",x"00",x"17", -- 0x13E8
    x"2E",x"45",x"5C",x"73",x"8A",x"A1",x"B8",x"CF", -- 0x13F0
    x"E6",x"FD",x"14",x"2B",x"42",x"59",x"70",x"87", -- 0x13F8
    x"9E",x"B5",x"CC",x"E3",x"FA",x"11",x"28",x"1E", -- 0x1400
    x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E", -- 0x1408
    x"1E",x"1E",x"1E",x"1F",x"1F",x"1F",x"1F",x"1F", -- 0x1410
    x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F", -- 0x1418
    x"1F",x"42",x"43",x"48",x"49",x"4E",x"4F",x"0B", -- 0x1420
    x"0A",x"09",x"08",x"07",x"06",x"05",x"04",x"03", -- 0x1428
    x"02",x"01",x"00",x"17",x"16",x"15",x"14",x"13", -- 0x1430
    x"12",x"11",x"10",x"0F",x"0E",x"0D",x"0C",x"23", -- 0x1438
    x"22",x"21",x"20",x"1F",x"1E",x"1D",x"1C",x"1B", -- 0x1440
    x"1A",x"19",x"18",x"2F",x"2E",x"2D",x"2C",x"2B", -- 0x1448
    x"2A",x"29",x"28",x"27",x"26",x"25",x"24",x"3B", -- 0x1450
    x"3A",x"39",x"38",x"37",x"36",x"35",x"34",x"33", -- 0x1458
    x"32",x"31",x"30",x"00",x"01",x"02",x"03",x"04", -- 0x1460
    x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C", -- 0x1468
    x"0D",x"0E",x"0F",x"10",x"11",x"12",x"13",x"14", -- 0x1470
    x"15",x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C", -- 0x1478
    x"1D",x"1E",x"1F",x"20",x"21",x"22",x"23",x"24", -- 0x1480
    x"25",x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C", -- 0x1488
    x"2D",x"2E",x"2F",x"30",x"31",x"32",x"33",x"34", -- 0x1490
    x"35",x"36",x"37",x"38",x"39",x"3A",x"3B",x"00", -- 0x1498
    x"00",x"00",x"00",x"00",x"40",x"30",x"20",x"10", -- 0x14A0
    x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x14A8
    x"01",x"01",x"01",x"01",x"00",x"00",x"01",x"01", -- 0x14B0
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x14B8
    x"00",x"00",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x14C0
    x"02",x"02",x"02",x"02",x"00",x"00",x"02",x"02", -- 0x14C8
    x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x14D0
    x"00",x"00",x"03",x"03",x"03",x"03",x"03",x"03", -- 0x14D8
    x"03",x"03",x"03",x"03",x"00",x"10",x"20",x"30", -- 0x14E0
    x"38",x"38",x"38",x"40",x"40",x"40",x"2E",x"5C", -- 0x14E8
    x"8A",x"A1",x"A1",x"A1",x"B8",x"B8",x"B8",x"1E", -- 0x14F0
    x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E", -- 0x14F8
    x"03",x"12",x"FF",x"02",x"07",x"07",x"7F",x"FF", -- 0x1500
    x"FF",x"FF",x"FF",x"13",x"F8",x"00",x"00",x"00", -- 0x1508
    x"F0",x"F8",x"F8",x"F8",x"F8",x"14",x"00",x"00", -- 0x1510
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02", -- 0x1518
    x"12",x"7F",x"01",x"03",x"03",x"3F",x"7F",x"7F", -- 0x1520
    x"7F",x"7F",x"13",x"FC",x"00",x"80",x"80",x"F8", -- 0x1528
    x"FC",x"FC",x"FC",x"FC",x"02",x"12",x"3F",x"00", -- 0x1530
    x"01",x"01",x"1F",x"3F",x"3F",x"3F",x"3F",x"13", -- 0x1538
    x"FE",x"80",x"C0",x"C0",x"FC",x"FE",x"FE",x"FE", -- 0x1540
    x"FE",x"03",x"12",x"1F",x"00",x"00",x"00",x"0F", -- 0x1548
    x"1F",x"1F",x"1F",x"1F",x"13",x"FF",x"40",x"E0", -- 0x1550
    x"E0",x"FE",x"FF",x"FF",x"FF",x"FF",x"14",x"00", -- 0x1558
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1560
    x"03",x"12",x"0F",x"00",x"00",x"00",x"07",x"0F", -- 0x1568
    x"0F",x"0F",x"0F",x"13",x"FF",x"20",x"70",x"70", -- 0x1570
    x"FF",x"FF",x"FF",x"FF",x"FF",x"14",x"80",x"00", -- 0x1578
    x"00",x"00",x"00",x"80",x"80",x"80",x"80",x"03", -- 0x1580
    x"12",x"07",x"00",x"00",x"00",x"03",x"07",x"07", -- 0x1588
    x"07",x"07",x"13",x"FF",x"10",x"38",x"38",x"FF", -- 0x1590
    x"FF",x"FF",x"FF",x"FF",x"14",x"C0",x"00",x"00", -- 0x1598
    x"00",x"80",x"C0",x"C0",x"C0",x"C0",x"03",x"12", -- 0x15A0
    x"03",x"00",x"00",x"00",x"01",x"03",x"03",x"03", -- 0x15A8
    x"03",x"13",x"FF",x"08",x"1C",x"1C",x"FF",x"FF", -- 0x15B0
    x"FF",x"FF",x"FF",x"14",x"E0",x"00",x"00",x"00", -- 0x15B8
    x"C0",x"E0",x"E0",x"E0",x"E0",x"03",x"12",x"01", -- 0x15C0
    x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01", -- 0x15C8
    x"13",x"FF",x"04",x"0E",x"0E",x"FF",x"FF",x"FF", -- 0x15D0
    x"FF",x"FF",x"14",x"F0",x"00",x"00",x"00",x"E0", -- 0x15D8
    x"F0",x"F0",x"F0",x"F0",x"89",x"22",x"7E",x"FF", -- 0x15E0
    x"FF",x"7E",x"24",x"91",x"00",x"00",x"00",x"00", -- 0x15E8
    x"00",x"00",x"00",x"00",x"44",x"11",x"3F",x"7F", -- 0x15F0
    x"7F",x"3F",x"12",x"48",x"80",x"00",x"00",x"80", -- 0x15F8
    x"80",x"00",x"00",x"80",x"22",x"08",x"1F",x"3F", -- 0x1600
    x"3F",x"1F",x"09",x"24",x"40",x"80",x"80",x"C0", -- 0x1608
    x"C0",x"80",x"00",x"40",x"11",x"04",x"0F",x"1F", -- 0x1610
    x"1F",x"0F",x"04",x"12",x"20",x"40",x"C0",x"E0", -- 0x1618
    x"E0",x"C0",x"80",x"20",x"08",x"02",x"07",x"0F", -- 0x1620
    x"0F",x"07",x"02",x"09",x"90",x"20",x"E0",x"F0", -- 0x1628
    x"F0",x"E0",x"40",x"10",x"04",x"01",x"03",x"07", -- 0x1630
    x"07",x"03",x"01",x"04",x"48",x"10",x"F0",x"F8", -- 0x1638
    x"F8",x"F0",x"20",x"88",x"02",x"00",x"01",x"03", -- 0x1640
    x"03",x"01",x"00",x"02",x"24",x"88",x"F8",x"FC", -- 0x1648
    x"FC",x"F8",x"90",x"44",x"01",x"00",x"00",x"01", -- 0x1650
    x"01",x"00",x"00",x"01",x"12",x"44",x"FC",x"FE", -- 0x1658
    x"FE",x"FC",x"48",x"22",x"38",x"78",x"BC",x"78", -- 0x1660
    x"B8",x"7C",x"B8",x"54",x"00",x"00",x"00",x"00", -- 0x1668
    x"00",x"00",x"00",x"00",x"0E",x"1E",x"2F",x"1E", -- 0x1670
    x"2E",x"1F",x"2E",x"15",x"00",x"00",x"00",x"00", -- 0x1678
    x"00",x"00",x"00",x"00",x"03",x"07",x"0B",x"07", -- 0x1680
    x"0B",x"07",x"0B",x"05",x"80",x"80",x"C0",x"80", -- 0x1688
    x"80",x"C0",x"80",x"40",x"00",x"01",x"02",x"01", -- 0x1690
    x"02",x"01",x"02",x"01",x"E0",x"E0",x"F0",x"E0", -- 0x1698
    x"E0",x"F0",x"E0",x"50",x"02",x"21",x"FD",x"08", -- 0x16A0
    x"45",x"20",x"10",x"C0",x"10",x"25",x"48",x"22", -- 0x16A8
    x"F8",x"80",x"10",x"20",x"40",x"18",x"40",x"20", -- 0x16B0
    x"90",x"02",x"21",x"3F",x"02",x"11",x"08",x"04", -- 0x16B8
    x"30",x"04",x"09",x"12",x"22",x"7E",x"20",x"44", -- 0x16C0
    x"08",x"10",x"06",x"10",x"48",x"24",x"02",x"21", -- 0x16C8
    x"0F",x"00",x"04",x"02",x"01",x"0C",x"01",x"02", -- 0x16D0
    x"04",x"22",x"DF",x"88",x"51",x"02",x"04",x"03", -- 0x16D8
    x"04",x"52",x"89",x"01",x"21",x"07",x"00",x"02", -- 0x16E0
    x"01",x"00",x"06",x"00",x"01",x"02",x"01",x"21", -- 0x16E8
    x"C7",x"00",x"82",x"C1",x"C0",x"C6",x"00",x"81", -- 0x16F0
    x"02",x"01",x"21",x"C7",x"00",x"02",x"01",x"80", -- 0x16F8
    x"C6",x"40",x"41",x"02",x"01",x"23",x"C0",x"00", -- 0x1700
    x"80",x"00",x"00",x"C0",x"00",x"00",x"80",x"01", -- 0x1708
    x"23",x"C3",x"00",x"81",x"03",x"03",x"C3",x"00", -- 0x1710
    x"01",x"80",x"01",x"23",x"C1",x"00",x"80",x"00", -- 0x1718
    x"00",x"C1",x"01",x"01",x"80",x"01",x"22",x"EF", -- 0x1720
    x"44",x"28",x"01",x"82",x"00",x"82",x"29",x"44", -- 0x1728
    x"64",x"63",x"00",x"64",x"80",x"64",x"63",x"7F", -- 0x1730
    x"80",x"41",x"7F",x"77",x"76",x"78",x"5A",x"78", -- 0x1738
    x"77",x"7F",x"80",x"5A",x"00",x"17",x"01",x"18", -- 0x1740
    x"0C",x"00",x"C0",x"30",x"85",x"CD",x"47",x"21", -- 0x1748
    x"68",x"63",x"DB",x"3A",x"62",x"E1",x"3B",x"9D", -- 0x1750
    x"03",x"4A",x"AD",x"A7",x"A5",x"A7",x"B0",x"A7", -- 0x1758
    x"AC",x"B0",x"B1",x"A3",x"A2",x"A2",x"A3",x"A3", -- 0x1760
    x"FF",x"FF",x"60",x"00",x"00",x"01",x"03",x"03", -- 0x1768
    x"03",x"03",x"03",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x1770
    x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x1778
    x"FF",x"FF",x"FF",x"00",x"00",x"80",x"C0",x"C0", -- 0x1780
    x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03", -- 0x1788
    x"03",x"03",x"03",x"FF",x"FF",x"FF",x"FF",x"F8", -- 0x1790
    x"F0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",x"1F", -- 0x1798
    x"0F",x"07",x"07",x"C0",x"C0",x"C0",x"C0",x"C0", -- 0x17A0
    x"C0",x"C0",x"C0",x"00",x"01",x"02",x"03",x"17", -- 0x17A8
    x"18",x"19",x"1A",x"05",x"06",x"07",x"08",x"1C", -- 0x17B0
    x"1D",x"1E",x"1F",x"0A",x"0B",x"0C",x"0D",x"21", -- 0x17B8
    x"22",x"23",x"24",x"0F",x"10",x"11",x"12",x"26", -- 0x17C0
    x"27",x"28",x"29",x"20",x"40",x"80",x"40",x"20", -- 0x17C8
    x"40",x"80",x"40",x"20",x"40",x"80",x"00",x"00", -- 0x17D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80", -- 0x17D8
    x"40",x"20",x"40",x"80",x"40",x"20",x"40",x"80", -- 0x17E0
    x"40",x"20",x"00",x"20",x"40",x"80",x"40",x"20", -- 0x17E8
    x"40",x"80",x"40",x"20",x"40",x"80",x"00",x"00", -- 0x17F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80", -- 0x17F8
    x"40",x"20",x"40",x"80",x"40",x"20",x"40",x"80", -- 0x1800
    x"40",x"20",x"00",x"08",x"10",x"20",x"10",x"08", -- 0x1808
    x"10",x"20",x"10",x"08",x"10",x"20",x"00",x"00", -- 0x1810
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20", -- 0x1818
    x"10",x"08",x"10",x"20",x"10",x"08",x"10",x"20", -- 0x1820
    x"10",x"08",x"00",x"08",x"10",x"20",x"10",x"08", -- 0x1828
    x"10",x"20",x"10",x"08",x"10",x"20",x"00",x"00", -- 0x1830
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20", -- 0x1838
    x"10",x"08",x"10",x"20",x"10",x"08",x"10",x"20", -- 0x1840
    x"10",x"08",x"00",x"02",x"04",x"08",x"04",x"02", -- 0x1848
    x"04",x"08",x"04",x"02",x"04",x"08",x"00",x"00", -- 0x1850
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08", -- 0x1858
    x"04",x"02",x"04",x"08",x"04",x"02",x"04",x"08", -- 0x1860
    x"04",x"02",x"00",x"02",x"04",x"08",x"04",x"02", -- 0x1868
    x"04",x"08",x"04",x"02",x"04",x"08",x"00",x"00", -- 0x1870
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08", -- 0x1878
    x"04",x"02",x"04",x"08",x"04",x"02",x"04",x"08", -- 0x1880
    x"04",x"02",x"00",x"40",x"40",x"40",x"40",x"40", -- 0x1888
    x"40",x"40",x"40",x"40",x"E0",x"40",x"00",x"00", -- 0x1890
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40", -- 0x1898
    x"40",x"40",x"40",x"40",x"40",x"E0",x"40",x"40", -- 0x18A0
    x"40",x"40",x"00",x"40",x"40",x"40",x"E0",x"40", -- 0x18A8
    x"40",x"40",x"40",x"40",x"40",x"40",x"00",x"00", -- 0x18B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0", -- 0x18B8
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x18C0
    x"40",x"40",x"00",x"10",x"10",x"10",x"10",x"10", -- 0x18C8
    x"10",x"10",x"10",x"10",x"38",x"10",x"00",x"00", -- 0x18D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10", -- 0x18D8
    x"10",x"10",x"10",x"10",x"10",x"38",x"10",x"10", -- 0x18E0
    x"10",x"10",x"00",x"10",x"10",x"10",x"38",x"10", -- 0x18E8
    x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00", -- 0x18F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38", -- 0x18F8
    x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10", -- 0x1900
    x"10",x"10",x"00",x"04",x"04",x"04",x"04",x"04", -- 0x1908
    x"04",x"04",x"04",x"04",x"0E",x"04",x"00",x"00", -- 0x1910
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04", -- 0x1918
    x"04",x"04",x"04",x"04",x"04",x"0E",x"04",x"04", -- 0x1920
    x"04",x"04",x"00",x"04",x"04",x"04",x"0E",x"04", -- 0x1928
    x"04",x"04",x"04",x"04",x"04",x"04",x"00",x"00", -- 0x1930
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1938
    x"0E",x"04",x"04",x"04",x"04",x"04",x"04",x"04", -- 0x1940
    x"04",x"04",x"00",x"40",x"40",x"40",x"40",x"40", -- 0x1948
    x"40",x"C0",x"60",x"C0",x"60",x"40",x"00",x"00", -- 0x1950
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40", -- 0x1958
    x"40",x"40",x"40",x"C0",x"60",x"C0",x"60",x"40", -- 0x1960
    x"40",x"40",x"00",x"40",x"40",x"C0",x"60",x"C0", -- 0x1968
    x"60",x"40",x"40",x"40",x"40",x"40",x"00",x"00", -- 0x1970
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0", -- 0x1978
    x"60",x"C0",x"60",x"40",x"40",x"40",x"40",x"40", -- 0x1980
    x"40",x"40",x"00",x"10",x"10",x"10",x"10",x"10", -- 0x1988
    x"10",x"30",x"18",x"30",x"18",x"10",x"00",x"00", -- 0x1990
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10", -- 0x1998
    x"10",x"10",x"10",x"18",x"30",x"18",x"30",x"10", -- 0x19A0
    x"10",x"10",x"00",x"10",x"10",x"30",x"18",x"30", -- 0x19A8
    x"18",x"10",x"10",x"10",x"10",x"10",x"00",x"00", -- 0x19B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- 0x19B8
    x"30",x"18",x"30",x"10",x"10",x"10",x"10",x"10", -- 0x19C0
    x"10",x"10",x"00",x"04",x"04",x"04",x"04",x"04", -- 0x19C8
    x"04",x"0C",x"06",x"0C",x"06",x"04",x"00",x"00", -- 0x19D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04", -- 0x19D8
    x"04",x"04",x"04",x"0C",x"06",x"0C",x"06",x"04", -- 0x19E0
    x"04",x"04",x"00",x"04",x"04",x"0C",x"06",x"0C", -- 0x19E8
    x"06",x"04",x"04",x"04",x"04",x"04",x"00",x"00", -- 0x19F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0C", -- 0x19F8
    x"06",x"0C",x"06",x"04",x"04",x"04",x"04",x"04", -- 0x1A00
    x"04",x"04",x"00",x"CB",x"8B",x"4B",x"B7",x"B8", -- 0x1A08
    x"B9",x"05",x"05",x"0A",x"08",x"0B",x"09",x"06", -- 0x1A10
    x"02",x"01",x"04",x"01",x"0B",x"09",x"09",x"0B", -- 0x1A18
    x"01",x"09",x"01",x"07",x"06",x"0A",x"01",x"09", -- 0x1A20
    x"04",x"0B",x"07",x"0A",x"06",x"01",x"06",x"01", -- 0x1A28
    x"06",x"06",x"0A",x"05",x"03",x"09",x"01",x"06", -- 0x1A30
    x"02",x"09",x"0A",x"07",x"01",x"01",x"02",x"0A", -- 0x1A38
    x"01",x"01",x"02",x"0B",x"06",x"0A",x"0B",x"0A", -- 0x1A40
    x"09",x"05",x"03",x"0B",x"05",x"08",x"01",x"0B", -- 0x1A48
    x"07",x"05",x"0B",x"05",x"01",x"08",x"0B",x"0B", -- 0x1A50
    x"01",x"07",x"02",x"06",x"01",x"0A",x"0B",x"04", -- 0x1A58
    x"02",x"01",x"09",x"0A",x"05",x"0A",x"0B",x"01", -- 0x1A60
    x"0B",x"0A",x"04",x"01",x"06",x"0B",x"01",x"08", -- 0x1A68
    x"01",x"02",x"0B",x"0A",x"0B",x"04",x"09",x"04", -- 0x1A70
    x"0A",x"0A",x"0B",x"0A",x"03",x"0B",x"01",x"09", -- 0x1A78
    x"0B",x"06",x"04",x"0A",x"06",x"04",x"02",x"02", -- 0x1A80
    x"09",x"0B",x"03",x"05",x"02",x"03",x"07",x"0B", -- 0x1A88
    x"02",x"05",x"0B",x"06",x"08",x"0B",x"08",x"01", -- 0x1A90
    x"0A",x"07",x"02",x"0B",x"01",x"01",x"06",x"08", -- 0x1A98
    x"01",x"08",x"09",x"0B",x"01",x"0B",x"0A",x"0B", -- 0x1AA0
    x"03",x"09",x"06",x"01",x"0A",x"0A",x"02",x"04", -- 0x1AA8
    x"0A",x"0B",x"09",x"02",x"07",x"08",x"04",x"01", -- 0x1AB0
    x"0B",x"06",x"02",x"0B",x"02",x"0A",x"0A",x"0B", -- 0x1AB8
    x"0B",x"08",x"07",x"0B",x"09",x"03",x"02",x"0B", -- 0x1AC0
    x"01",x"0B",x"01",x"05",x"01",x"01",x"06",x"03", -- 0x1AC8
    x"04",x"03",x"02",x"0B",x"0B",x"08",x"01",x"0B", -- 0x1AD0
    x"01",x"06",x"0A",x"03",x"08",x"01",x"0A",x"02", -- 0x1AD8
    x"07",x"07",x"06",x"01",x"05",x"05",x"09",x"01", -- 0x1AE0
    x"01",x"07",x"07",x"0B",x"0A",x"04",x"08",x"01", -- 0x1AE8
    x"01",x"07",x"0B",x"02",x"0B",x"0A",x"0A",x"08", -- 0x1AF0
    x"06",x"02",x"08",x"06",x"0B",x"01",x"06",x"0A", -- 0x1AF8
    x"0B",x"09",x"0B",x"07",x"02",x"0A",x"0B",x"02", -- 0x1B00
    x"07",x"0B",x"02",x"0B",x"0B",x"01",x"04",x"08", -- 0x1B08
    x"0A",x"03",x"25",x"FF",x"03",x"0F",x"1F",x"3F", -- 0x1B10
    x"6D",x"FF",x"38",x"10",x"26",x"FF",x"C0",x"F0", -- 0x1B18
    x"F8",x"FC",x"B6",x"FF",x"1C",x"08",x"27",x"00", -- 0x1B20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B28
    x"03",x"25",x"3F",x"00",x"03",x"07",x"0F",x"1B", -- 0x1B30
    x"3F",x"0E",x"04",x"26",x"FF",x"F0",x"FC",x"FE", -- 0x1B38
    x"FF",x"6D",x"FF",x"07",x"02",x"27",x"C0",x"00", -- 0x1B40
    x"00",x"00",x"00",x"80",x"C0",x"00",x"00",x"03", -- 0x1B48
    x"25",x"0F",x"00",x"00",x"01",x"03",x"06",x"0F", -- 0x1B50
    x"03",x"01",x"26",x"FF",x"3C",x"FF",x"FF",x"FF", -- 0x1B58
    x"DB",x"FF",x"81",x"00",x"27",x"F0",x"00",x"00", -- 0x1B60
    x"80",x"C0",x"60",x"F0",x"C0",x"80",x"03",x"25", -- 0x1B68
    x"03",x"00",x"00",x"00",x"00",x"01",x"03",x"00", -- 0x1B70
    x"00",x"26",x"FF",x"0F",x"3F",x"7F",x"FF",x"B6", -- 0x1B78
    x"FF",x"E0",x"40",x"27",x"FC",x"00",x"C0",x"E0", -- 0x1B80
    x"F0",x"D8",x"FC",x"70",x"20",x"03",x"25",x"BF", -- 0x1B88
    x"25",x"10",x"A3",x"07",x"0F",x"27",x"83",x"1E", -- 0x1B90
    x"26",x"FF",x"22",x"08",x"C4",x"F2",x"EA",x"E0", -- 0x1B98
    x"60",x"1E",x"27",x"80",x"00",x"00",x"80",x"00", -- 0x1BA0
    x"00",x"00",x"80",x"00",x"03",x"25",x"2F",x"09", -- 0x1BA8
    x"04",x"28",x"01",x"03",x"09",x"20",x"08",x"26", -- 0x1BB0
    x"FF",x"48",x"02",x"F1",x"FC",x"FA",x"F8",x"D8", -- 0x1BB8
    x"80",x"27",x"E0",x"80",x"00",x"20",x"80",x"80", -- 0x1BC0
    x"00",x"20",x"20",x"03",x"25",x"0B",x"02",x"01", -- 0x1BC8
    x"0A",x"00",x"00",x"02",x"08",x"00",x"26",x"FF", -- 0x1BD0
    x"52",x"00",x"3C",x"7F",x"FE",x"7E",x"36",x"10", -- 0x1BD8
    x"27",x"F8",x"20",x"80",x"48",x"20",x"A0",x"00", -- 0x1BE0
    x"08",x"50",x"03",x"25",x"02",x"00",x"00",x"02", -- 0x1BE8
    x"00",x"00",x"00",x"02",x"00",x"26",x"FF",x"94", -- 0x1BF0
    x"40",x"8F",x"1F",x"3F",x"9F",x"0D",x"80",x"27", -- 0x1BF8
    x"FE",x"88",x"20",x"12",x"C8",x"A8",x"80",x"82", -- 0x1C00
    x"60",x"30",x"05",x"10",x"10",x"15",x"10",x"05", -- 0x1C08
    x"05",x"10",x"10",x"15",x"05",x"05",x"10",x"10", -- 0x1C10
    x"03",x"12",x"BF",x"0A",x"82",x"0A",x"02",x"82", -- 0x1C18
    x"A6",x"1F",x"3F",x"13",x"FF",x"02",x"0C",x"70", -- 0x1C20
    x"02",x"18",x"C0",x"F9",x"F9",x"14",x"80",x"00", -- 0x1C28
    x"00",x"80",x"00",x"80",x"00",x"00",x"80",x"03", -- 0x1C30
    x"12",x"2F",x"02",x"20",x"02",x"00",x"20",x"29", -- 0x1C38
    x"07",x"0F",x"13",x"FF",x"80",x"83",x"9C",x"80", -- 0x1C40
    x"86",x"B0",x"FE",x"FE",x"14",x"E0",x"80",x"00", -- 0x1C48
    x"20",x"80",x"20",x"00",x"40",x"60",x"03",x"12", -- 0x1C50
    x"0B",x"00",x"08",x"00",x"00",x"08",x"0A",x"01", -- 0x1C58
    x"03",x"13",x"FF",x"A0",x"20",x"A7",x"20",x"21", -- 0x1C60
    x"6C",x"FF",x"FF",x"14",x"F8",x"20",x"C0",x"08", -- 0x1C68
    x"20",x"88",x"00",x"90",x"98",x"03",x"12",x"02", -- 0x1C70
    x"00",x"02",x"00",x"00",x"02",x"02",x"00",x"00", -- 0x1C78
    x"13",x"FF",x"28",x"08",x"29",x"08",x"08",x"9B", -- 0x1C80
    x"7F",x"FF",x"14",x"FE",x"08",x"30",x"C2",x"08", -- 0x1C88
    x"62",x"00",x"E4",x"E6",x"03",x"12",x"FF",x"03", -- 0x1C90
    x"40",x"04",x"A0",x"09",x"42",x"1F",x"3F",x"13", -- 0x1C98
    x"FF",x"08",x"40",x"14",x"81",x"25",x"00",x"F4", -- 0x1CA0
    x"F7",x"14",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA8
    x"00",x"00",x"00",x"03",x"12",x"3F",x"00",x"10", -- 0x1CB0
    x"01",x"28",x"02",x"10",x"07",x"0F",x"13",x"FF", -- 0x1CB8
    x"C2",x"10",x"05",x"20",x"49",x"80",x"FD",x"FD", -- 0x1CC0
    x"14",x"C0",x"00",x"00",x"00",x"40",x"40",x"00", -- 0x1CC8
    x"00",x"C0",x"03",x"12",x"0F",x"00",x"04",x"00", -- 0x1CD0
    x"0A",x"00",x"04",x"01",x"03",x"13",x"FF",x"30", -- 0x1CD8
    x"04",x"41",x"08",x"92",x"20",x"FF",x"FF",x"14", -- 0x1CE0
    x"F0",x"80",x"00",x"40",x"10",x"50",x"00",x"40", -- 0x1CE8
    x"70",x"03",x"12",x"03",x"00",x"01",x"00",x"02", -- 0x1CF0
    x"00",x"01",x"00",x"00",x"13",x"FF",x"20",x"02", -- 0x1CF8
    x"10",x"44",x"21",x"02",x"7F",x"FF",x"14",x"FF", -- 0x1D00
    x"88",x"22",x"00",x"81",x"12",x"00",x"D0",x"DC", -- 0x1D08
    x"01",x"14",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D10
    x"00",x"00",x"00",x"07",x"01",x"0D",x"05",x"20", -- 0x1D18
    x"0F",x"16",x"05",x"12",x"F0",x"09",x"02",x"20", -- 0x1D20
    x"20",x"20",x"20",x"F0",x"05",x"04",x"09",x"0E", -- 0x1D28
    x"13",x"14",x"12",x"15",x"03",x"14",x"09",x"0F", -- 0x1D30
    x"0E",x"13",x"F0",x"00",x"06",x"FE",x"00",x"2A", -- 0x1D38
    x"20",x"13",x"03",x"0F",x"12",x"05",x"20",x"01", -- 0x1D40
    x"04",x"16",x"01",x"0E",x"03",x"05",x"20",x"14", -- 0x1D48
    x"01",x"02",x"0C",x"05",x"20",x"2A",x"F0",x"05", -- 0x1D50
    x"08",x"65",x"66",x"67",x"F0",x"05",x"0A",x"4E", -- 0x1D58
    x"4F",x"F0",x"05",x"0C",x"48",x"49",x"F0",x"05", -- 0x1D60
    x"0E",x"42",x"43",x"F0",x"08",x"08",x"FE",x"0A", -- 0x1D68
    x"3D",x"3F",x"20",x"0D",x"19",x"13",x"14",x"05", -- 0x1D70
    x"12",x"19",x"F0",x"08",x"0A",x"3D",x"33",x"30", -- 0x1D78
    x"20",x"10",x"0F",x"09",x"0E",x"14",x"13",x"F0", -- 0x1D80
    x"08",x"0C",x"3D",x"32",x"30",x"20",x"10",x"0F", -- 0x1D88
    x"09",x"0E",x"14",x"13",x"F0",x"08",x"0E",x"3D", -- 0x1D90
    x"31",x"30",x"20",x"10",x"0F",x"09",x"0E",x"14", -- 0x1D98
    x"13",x"F0",x"01",x"10",x"15",x"13",x"05",x"20", -- 0x1DA0
    x"0A",x"0F",x"19",x"13",x"14",x"09",x"03",x"0B", -- 0x1DA8
    x"20",x"0F",x"12",x"20",x"0B",x"05",x"19",x"13", -- 0x1DB0
    x"2E",x"F0",x"01",x"12",x"8C",x"2D",x"0C",x"05", -- 0x1DB8
    x"06",x"14",x"20",x"8D",x"2D",x"06",x"09",x"12", -- 0x1DC0
    x"05",x"20",x"8E",x"2D",x"12",x"09",x"07",x"08", -- 0x1DC8
    x"14",x"F0",x"00",x"14",x"14",x"0F",x"10",x"20", -- 0x1DD0
    x"31",x"35",x"30",x"30",x"20",x"06",x"0F",x"12", -- 0x1DD8
    x"20",x"05",x"18",x"14",x"12",x"01",x"20",x"02", -- 0x1DE0
    x"01",x"13",x"05",x"FE",x"78",x"20",x"FF",x"E5", -- 0x1DE8
    x"E1",x"DF",x"DD",x"00",x"F7",x"ED",x"E2",x"D8", -- 0x1DF0
    x"00",x"00",x"BD",x"C7",x"D2",x"DC",x"E6",x"00", -- 0x1DF8
    x"FB",x"F9",x"00",x"F3",x"00",x"E8",x"00",x"D0", -- 0x1E00
    x"F5",x"F6",x"F7",x"F8",x"F9",x"F8",x"F7",x"F6", -- 0x1E08
    x"F5",x"F4",x"F3",x"F2",x"01",x"04",x"05",x"05", -- 0x1E10
    x"06",x"06",x"06",x"06",x"04",x"04",x"04",x"04", -- 0x1E18
    x"07",x"07",x"07",x"07",x"07",x"02",x"02",x"02", -- 0x1E20
    x"03",x"03",x"13",x"03",x"30",x"30",x"30",x"30", -- 0x1E28
    x"30",x"20",x"08",x"09",x"30",x"30",x"30",x"30", -- 0x1E30
    x"30",x"20",x"30",x"7C",x"42",x"42",x"7C",x"40", -- 0x1E38
    x"40",x"40",x"00",x"42",x"42",x"42",x"42",x"42", -- 0x1E40
    x"42",x"3C",x"00",x"3C",x"42",x"40",x"3C",x"02", -- 0x1E48
    x"42",x"3C",x"00",x"42",x"42",x"42",x"7E",x"42", -- 0x1E50
    x"42",x"42",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E58
    x"00",x"00",x"00",x"F2",x"86",x"82",x"E2",x"82", -- 0x1E60
    x"82",x"87",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E68
    x"00",x"00",x"00",x"3E",x"08",x"08",x"08",x"08", -- 0x1E70
    x"08",x"08",x"00",x"18",x"24",x"42",x"42",x"42", -- 0x1E78
    x"24",x"18",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E80
    x"00",x"00",x"00",x"7C",x"22",x"22",x"3C",x"22", -- 0x1E88
    x"22",x"7C",x"00",x"7E",x"40",x"40",x"78",x"40", -- 0x1E90
    x"40",x"7E",x"00",x"1C",x"22",x"40",x"4E",x"42", -- 0x1E98
    x"22",x"1C",x"00",x"1C",x"08",x"08",x"08",x"08", -- 0x1EA0
    x"08",x"1C",x"00",x"42",x"62",x"52",x"4A",x"46", -- 0x1EA8
    x"42",x"42",x"00",x"A5",x"A5",x"A5",x"BD",x"81", -- 0x1EB0
    x"BD",x"A5",x"E5",x"18",x"24",x"24",x"5A",x"42", -- 0x1EB8
    x"99",x"A5",x"A5",x"E0",x"A0",x"A0",x"A0",x"A0", -- 0x1EC0
    x"BF",x"81",x"BF",x"00",x"00",x"00",x"00",x"00", -- 0x1EC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED0
    x"00",x"00",x"00",x"7E",x"BD",x"81",x"BC",x"7E", -- 0x1ED8
    x"01",x"BD",x"7E",x"00",x"00",x"00",x"00",x"00", -- 0x1EE0
    x"38",x"28",x"28",x"C3",x"A5",x"99",x"A5",x"BD", -- 0x1EE8
    x"A5",x"A5",x"E5",x"18",x"24",x"24",x"5A",x"42", -- 0x1EF0
    x"99",x"A5",x"A5",x"FE",x"82",x"EE",x"28",x"28", -- 0x1EF8
    x"28",x"28",x"28",x"7E",x"BD",x"81",x"BC",x"7E", -- 0x1F00
    x"01",x"BD",x"7E",x"55",x"55",x"55",x"55",x"55", -- 0x1F08
    x"5D",x"41",x"3E",x"3E",x"41",x"5D",x"55",x"55", -- 0x1F10
    x"5D",x"41",x"3E",x"53",x"55",x"5A",x"54",x"44", -- 0x1F18
    x"52",x"59",x"77",x"18",x"24",x"24",x"5A",x"42", -- 0x1F20
    x"99",x"A5",x"A5",x"10",x"0C",x"01",x"19",x"20", -- 0x1F28
    x"10",x"0C",x"01",x"19",x"05",x"12",x"20",x"31", -- 0x1F30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"30", -- 0x1F38
    x"99",x"A5",x"A5",x"E0",x"A0",x"A0",x"A0",x"A0", -- 0x1F40
    x"BF",x"81",x"BF",x"00",x"00",x"00",x"00",x"00", -- 0x1F48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F50
    x"00",x"00",x"00",x"7E",x"BD",x"81",x"BC",x"7E", -- 0x1F58
    x"01",x"BD",x"7E",x"00",x"00",x"00",x"00",x"00", -- 0x1F60
    x"38",x"28",x"28",x"C3",x"A5",x"99",x"A5",x"BD", -- 0x1F68
    x"A5",x"A5",x"E5",x"18",x"24",x"24",x"5A",x"42", -- 0x1F70
    x"99",x"A5",x"A5",x"FE",x"00",x"43",x"C0",x"2B", -- 0x1F78
    x"03",x"47",x"65",x"73",x"B5",x"A1",x"FC",x"93", -- 0x1F80
    x"20",x"D3",x"49",x"5A",x"C6",x"13",x"D3",x"D3", -- 0x1F88
    x"35",x"89",x"05",x"2C",x"3D",x"18",x"78",x"F2", -- 0x1F90
    x"80",x"C2",x"08",x"95",x"09",x"42",x"44",x"12", -- 0x1F98
    x"8D",x"C5",x"D4",x"8B",x"7C",x"5E",x"BC",x"7F", -- 0x1FA0
    x"3F",x"95",x"E8",x"6D",x"0C",x"0C",x"8C",x"38", -- 0x1FA8
    x"9E",x"09",x"8D",x"E2",x"34",x"FE",x"6E",x"3F", -- 0x1FB0
    x"78",x"76",x"0C",x"78",x"37",x"12",x"08",x"43", -- 0x1FB8
    x"25",x"4B",x"08",x"A2",x"1A",x"B3",x"F5",x"41", -- 0x1FC0
    x"A6",x"F7",x"90",x"DB",x"F3",x"C3",x"85",x"71", -- 0x1FC8
    x"6E",x"01",x"59",x"A2",x"3A",x"D0",x"8F",x"0B", -- 0x1FD0
    x"E0",x"E0",x"D7",x"E6",x"0C",x"0A",x"86",x"81", -- 0x1FD8
    x"EA",x"44",x"7E",x"6D",x"F4",x"DF",x"5C",x"03", -- 0x1FE0
    x"8C",x"FC",x"38",x"B3",x"2C",x"9F",x"A4",x"84", -- 0x1FE8
    x"6C",x"93",x"84",x"93",x"CC",x"16",x"5D",x"CF", -- 0x1FF0
    x"B8",x"32",x"FC",x"FB",x"9C",x"B3",x"25",x"23"  -- 0x1FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
