-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity cart_rom is --4K
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of cart_rom is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"09",x"A0",x"09",x"A0",x"41",x"30",x"C3",x"C2", -- 0x0000
    x"CD",x"4C",x"00",x"AF",x"78",x"D8",x"A9",x"00", -- 0x0008
    x"8D",x"21",x"02",x"8D",x"22",x"02",x"20",x"25", -- 0x0010
    x"19",x"A2",x"FF",x"9A",x"20",x"21",x"17",x"20", -- 0x0018
    x"17",x"18",x"20",x"6F",x"1A",x"20",x"97",x"10", -- 0x0020
    x"20",x"0D",x"11",x"20",x"5B",x"19",x"20",x"3E", -- 0x0028
    x"12",x"20",x"E6",x"12",x"20",x"CF",x"15",x"20", -- 0x0030
    x"7A",x"18",x"4C",x"1F",x"10",x"A0",x"0F",x"B9", -- 0x0038
    x"EA",x"13",x"99",x"00",x"90",x"88",x"10",x"F7", -- 0x0040
    x"60",x"A2",x"08",x"BD",x"30",x"14",x"95",x"20", -- 0x0048
    x"95",x"40",x"CA",x"10",x"F6",x"AE",x"23",x"02", -- 0x0050
    x"BD",x"A1",x"1B",x"85",x"23",x"85",x"43",x"60", -- 0x0058
    x"A2",x"00",x"A9",x"07",x"A0",x"05",x"18",x"95", -- 0x0060
    x"60",x"94",x"9D",x"69",x"08",x"E8",x"E0",x"08", -- 0x0068
    x"D0",x"F4",x"A2",x"04",x"18",x"A5",x"52",x"69", -- 0x0070
    x"09",x"A8",x"94",x"68",x"88",x"88",x"CA",x"10", -- 0x0078
    x"F9",x"A2",x"27",x"A9",x"01",x"95",x"6D",x"CA", -- 0x0080
    x"10",x"FB",x"A9",x"FF",x"85",x"9B",x"A9",x"09", -- 0x0088
    x"85",x"0B",x"85",x"0E",x"85",x"C2",x"60",x"C6", -- 0x0090
    x"20",x"D0",x"4D",x"A5",x"40",x"85",x"20",x"A5", -- 0x0098
    x"10",x"30",x"46",x"F0",x"43",x"A5",x"02",x"30", -- 0x00A0
    x"19",x"F0",x"26",x"A6",x"00",x"E0",x"50",x"F0", -- 0x00A8
    x"20",x"E8",x"86",x"01",x"A5",x"00",x"20",x"2B", -- 0x00B0
    x"12",x"AD",x"BB",x"13",x"99",x"A4",x"1F",x"4C", -- 0x00B8
    x"D1",x"10",x"A6",x"00",x"F0",x"0B",x"CA",x"86", -- 0x00C0
    x"01",x"A5",x"00",x"20",x"2B",x"12",x"C8",x"D0", -- 0x00C8
    x"E8",x"A5",x"01",x"85",x"00",x"20",x"2B",x"12", -- 0x00D0
    x"20",x"32",x"12",x"BD",x"BC",x"13",x"99",x"A4", -- 0x00D8
    x"1F",x"C8",x"BD",x"C0",x"13",x"99",x"A4",x"1F", -- 0x00E0
    x"60",x"C9",x"80",x"D0",x"13",x"A5",x"00",x"20", -- 0x00E8
    x"2B",x"12",x"AD",x"BB",x"13",x"99",x"A4",x"1F", -- 0x00F0
    x"C8",x"99",x"A4",x"1F",x"A9",x"01",x"85",x"C6", -- 0x00F8
    x"E6",x"10",x"A5",x"10",x"C9",x"A0",x"D0",x"04", -- 0x0100
    x"A9",x"00",x"85",x"10",x"60",x"C6",x"21",x"D0", -- 0x0108
    x"33",x"A5",x"41",x"85",x"21",x"A5",x"11",x"F0", -- 0x0110
    x"2B",x"30",x"29",x"C9",x"01",x"D0",x"26",x"A5", -- 0x0118
    x"10",x"30",x"21",x"F0",x"1F",x"18",x"A5",x"00", -- 0x0120
    x"69",x"02",x"85",x"03",x"20",x"2B",x"12",x"84", -- 0x0128
    x"05",x"20",x"32",x"12",x"86",x"06",x"A9",x"9F", -- 0x0130
    x"85",x"04",x"A9",x"02",x"85",x"11",x"20",x"F5", -- 0x0138
    x"11",x"4C",x"6B",x"11",x"60",x"A5",x"09",x"D0", -- 0x0140
    x"28",x"20",x"F5",x"11",x"A4",x"05",x"B1",x"07", -- 0x0148
    x"38",x"C9",x"2E",x"90",x"07",x"C9",x"3E",x"B0", -- 0x0150
    x"03",x"4C",x"63",x"11",x"A4",x"05",x"AD",x"BB", -- 0x0158
    x"13",x"91",x"07",x"C6",x"04",x"A5",x"04",x"C9", -- 0x0160
    x"FF",x"F0",x"2F",x"20",x"EB",x"11",x"4C",x"79", -- 0x0168
    x"11",x"C6",x"04",x"A5",x"04",x"18",x"4A",x"4A", -- 0x0170
    x"4A",x"85",x"0C",x"A4",x"04",x"20",x"10",x"12", -- 0x0178
    x"85",x"09",x"20",x"1A",x"12",x"20",x"39",x"14", -- 0x0180
    x"20",x"FD",x"18",x"A4",x"05",x"B1",x"07",x"4C", -- 0x0188
    x"9F",x"11",x"A4",x"05",x"AD",x"E9",x"13",x"91", -- 0x0190
    x"07",x"60",x"A9",x"80",x"85",x"11",x"60",x"38", -- 0x0198
    x"C9",x"2E",x"90",x"EE",x"C9",x"3E",x"B0",x"EA", -- 0x01A0
    x"85",x"56",x"38",x"E9",x"2E",x"85",x"57",x"0A", -- 0x01A8
    x"0A",x"0A",x"18",x"65",x"09",x"85",x"58",x"A8", -- 0x01B0
    x"B9",x"70",x"1D",x"A4",x"06",x"39",x"28",x"14", -- 0x01B8
    x"D0",x"07",x"A5",x"56",x"A4",x"05",x"91",x"07", -- 0x01C0
    x"60",x"B9",x"2C",x"14",x"85",x"5A",x"A5",x"58", -- 0x01C8
    x"A8",x"38",x"E9",x"02",x"85",x"5B",x"B9",x"70", -- 0x01D0
    x"1D",x"25",x"5A",x"99",x"70",x"1D",x"88",x"C4", -- 0x01D8
    x"5B",x"D0",x"F3",x"A9",x"80",x"85",x"11",x"4C", -- 0x01E0
    x"C2",x"11",x"60",x"A5",x"04",x"20",x"00",x"12", -- 0x01E8
    x"86",x"07",x"84",x"08",x"60",x"A0",x"07",x"A9", -- 0x01F0
    x"00",x"99",x"F0",x"1D",x"88",x"10",x"FA",x"60", -- 0x01F8
    x"18",x"4A",x"4A",x"4A",x"48",x"A8",x"B9",x"FA", -- 0x0200
    x"13",x"AA",x"B9",x"11",x"14",x"A8",x"68",x"60", -- 0x0208
    x"0A",x"0A",x"0A",x"85",x"F0",x"38",x"98",x"E5", -- 0x0210
    x"F0",x"60",x"A4",x"09",x"A6",x"06",x"BD",x"28", -- 0x0218
    x"14",x"99",x"F0",x"1D",x"C8",x"A9",x"00",x"99", -- 0x0220
    x"F0",x"1D",x"60",x"48",x"18",x"4A",x"4A",x"A8", -- 0x0228
    x"68",x"60",x"48",x"98",x"0A",x"0A",x"85",x"F0", -- 0x0230
    x"38",x"68",x"E5",x"F0",x"AA",x"60",x"C6",x"23", -- 0x0238
    x"D0",x"78",x"A5",x"43",x"85",x"23",x"C6",x"0B", -- 0x0240
    x"D0",x"70",x"A5",x"0E",x"85",x"0B",x"20",x"BB", -- 0x0248
    x"12",x"A9",x"10",x"85",x"C5",x"A5",x"9C",x"D0", -- 0x0250
    x"33",x"A5",x"9B",x"30",x"15",x"A5",x"96",x"C9", -- 0x0258
    x"03",x"D0",x"07",x"A9",x"AC",x"A2",x"13",x"20", -- 0x0260
    x"A7",x"12",x"A9",x"F6",x"8D",x"84",x"12",x"4C", -- 0x0268
    x"82",x"12",x"A5",x"96",x"D0",x"07",x"A9",x"A3", -- 0x0270
    x"A2",x"13",x"20",x"A7",x"12",x"A9",x"D6",x"8D", -- 0x0278
    x"84",x"12",x"A2",x"07",x"F6",x"60",x"CA",x"10", -- 0x0280
    x"FB",x"4C",x"EE",x"12",x"A9",x"B4",x"A2",x"13", -- 0x0288
    x"20",x"A7",x"12",x"A2",x"04",x"F6",x"68",x"CA", -- 0x0290
    x"10",x"FB",x"A5",x"9B",x"49",x"FE",x"85",x"9B", -- 0x0298
    x"A9",x"00",x"85",x"9C",x"4C",x"EE",x"12",x"8D", -- 0x02A0
    x"38",x"13",x"8E",x"39",x"13",x"20",x"EE",x"12", -- 0x02A8
    x"A9",x"72",x"8D",x"38",x"13",x"A9",x"13",x"8D", -- 0x02B0
    x"39",x"13",x"60",x"A5",x"9B",x"30",x"0F",x"A2", -- 0x02B8
    x"07",x"B5",x"9D",x"D0",x"1A",x"CA",x"10",x"F9", -- 0x02C0
    x"60",x"B5",x"60",x"F0",x"0D",x"60",x"A2",x"00", -- 0x02C8
    x"B5",x"9D",x"D0",x"F5",x"E8",x"E0",x"08",x"D0", -- 0x02D0
    x"F7",x"60",x"A9",x"01",x"85",x"9C",x"60",x"B5", -- 0x02D8
    x"60",x"C9",x"50",x"F0",x"F5",x"60",x"C6",x"24", -- 0x02E0
    x"D0",x"69",x"A5",x"44",x"85",x"24",x"A2",x"00", -- 0x02E8
    x"B5",x"9D",x"D0",x"06",x"E8",x"E0",x"08",x"D0", -- 0x02F0
    x"F7",x"60",x"86",x"0D",x"B5",x"60",x"20",x"2B", -- 0x02F8
    x"12",x"84",x"95",x"84",x"9A",x"20",x"32",x"12", -- 0x0300
    x"85",x"96",x"A2",x"00",x"86",x"97",x"A5",x"0D", -- 0x0308
    x"85",x"98",x"A5",x"95",x"85",x"9A",x"A6",x"97", -- 0x0310
    x"B4",x"68",x"B9",x"FA",x"13",x"8D",x"9B",x"13", -- 0x0318
    x"8D",x"A0",x"13",x"B9",x"11",x"14",x"8D",x"9C", -- 0x0320
    x"13",x"8D",x"A1",x"13",x"20",x"54",x"13",x"A6", -- 0x0328
    x"99",x"B5",x"6D",x"F0",x"05",x"30",x"29",x"20", -- 0x0330
    x"72",x"13",x"E6",x"99",x"18",x"A5",x"9A",x"69", -- 0x0338
    x"02",x"85",x"9A",x"E6",x"98",x"A5",x"98",x"C9", -- 0x0340
    x"08",x"D0",x"E4",x"E6",x"97",x"A5",x"97",x"C9", -- 0x0348
    x"05",x"D0",x"BB",x"60",x"18",x"A5",x"97",x"0A", -- 0x0350
    x"0A",x"0A",x"18",x"65",x"98",x"85",x"99",x"60", -- 0x0358
    x"A9",x"00",x"95",x"6D",x"AD",x"BB",x"13",x"AA", -- 0x0360
    x"20",x"98",x"13",x"A6",x"98",x"D6",x"9D",x"4C", -- 0x0368
    x"3A",x"13",x"A4",x"96",x"A5",x"97",x"F0",x"19", -- 0x0370
    x"38",x"C9",x"03",x"90",x"0A",x"B9",x"C8",x"13", -- 0x0378
    x"AA",x"B9",x"C4",x"13",x"4C",x"98",x"13",x"B9", -- 0x0380
    x"D0",x"13",x"AA",x"B9",x"CC",x"13",x"4C",x"98", -- 0x0388
    x"13",x"B9",x"D8",x"13",x"AA",x"B9",x"D4",x"13", -- 0x0390
    x"A4",x"9A",x"99",x"FF",x"FF",x"8A",x"C8",x"99", -- 0x0398
    x"FF",x"FF",x"60",x"A4",x"9A",x"AD",x"BB",x"13", -- 0x03A0
    x"C8",x"4C",x"9F",x"13",x"A4",x"9A",x"AD",x"BB", -- 0x03A8
    x"13",x"4C",x"9F",x"13",x"AD",x"BB",x"13",x"AA", -- 0x03B0
    x"4C",x"98",x"13",x"00",x"01",x"02",x"03",x"04", -- 0x03B8
    x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C", -- 0x03C0
    x"0D",x"0E",x"0F",x"10",x"11",x"12",x"13",x"14", -- 0x03C8
    x"15",x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C", -- 0x03D0
    x"1D",x"1E",x"1F",x"20",x"21",x"22",x"23",x"24", -- 0x03D8
    x"25",x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C", -- 0x03E0
    x"2D",x"3E",x"06",x"19",x"95",x"2E",x"00",x"FF", -- 0x03E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F0
    x"0F",x"6F",x"00",x"15",x"2A",x"3F",x"54",x"69", -- 0x03F8
    x"7E",x"93",x"A8",x"BD",x"D2",x"E7",x"FC",x"11", -- 0x0400
    x"26",x"3B",x"50",x"65",x"7A",x"8F",x"A4",x"B9", -- 0x0408
    x"CE",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E", -- 0x0410
    x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1F",x"1F", -- 0x0418
    x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F", -- 0x0420
    x"80",x"20",x"08",x"02",x"3F",x"CF",x"F3",x"FC", -- 0x0428
    x"70",x"0C",x"80",x"90",x"20",x"2A",x"D0",x"80", -- 0x0430
    x"09",x"A2",x"04",x"B5",x"68",x"C5",x"0C",x"F0", -- 0x0438
    x"04",x"CA",x"10",x"F7",x"60",x"8A",x"85",x"A9", -- 0x0440
    x"0A",x"0A",x"0A",x"85",x"A5",x"A2",x"07",x"38", -- 0x0448
    x"B5",x"60",x"C5",x"03",x"B0",x"34",x"69",x"04", -- 0x0450
    x"38",x"C5",x"03",x"90",x"2D",x"18",x"8A",x"65", -- 0x0458
    x"A5",x"A8",x"B9",x"6D",x"00",x"F0",x"DD",x"A9", -- 0x0460
    x"80",x"99",x"6D",x"00",x"85",x"11",x"A6",x"A9", -- 0x0468
    x"BD",x"0C",x"1B",x"20",x"8E",x"14",x"A5",x"43", -- 0x0470
    x"38",x"C9",x"09",x"90",x"08",x"AE",x"23",x"02", -- 0x0478
    x"FD",x"AB",x"1B",x"85",x"43",x"A9",x"01",x"85", -- 0x0480
    x"C6",x"60",x"CA",x"10",x"C2",x"60",x"F8",x"18", -- 0x0488
    x"6D",x"21",x"02",x"8D",x"21",x"02",x"90",x"08", -- 0x0490
    x"A9",x"00",x"6D",x"22",x"02",x"8D",x"22",x"02", -- 0x0498
    x"D8",x"A5",x"51",x"D0",x"0C",x"AD",x"22",x"02", -- 0x04A0
    x"F0",x"07",x"85",x"51",x"E6",x"50",x"20",x"3E", -- 0x04A8
    x"15",x"20",x"20",x"15",x"AD",x"22",x"02",x"20", -- 0x04B0
    x"18",x"15",x"A0",x"00",x"20",x"E2",x"14",x"AD", -- 0x04B8
    x"22",x"02",x"29",x"0F",x"A0",x"08",x"20",x"E2", -- 0x04C0
    x"14",x"AD",x"21",x"02",x"20",x"18",x"15",x"A0", -- 0x04C8
    x"10",x"20",x"E2",x"14",x"AD",x"21",x"02",x"29", -- 0x04D0
    x"0F",x"A0",x"18",x"20",x"E2",x"14",x"A9",x"00", -- 0x04D8
    x"A0",x"20",x"AA",x"A5",x"13",x"D0",x"49",x"BD", -- 0x04E0
    x"11",x"1B",x"99",x"48",x"1D",x"BD",x"1B",x"1B", -- 0x04E8
    x"99",x"49",x"1D",x"BD",x"25",x"1B",x"99",x"4A", -- 0x04F0
    x"1D",x"BD",x"2F",x"1B",x"99",x"4B",x"1D",x"BD", -- 0x04F8
    x"39",x"1B",x"99",x"4C",x"1D",x"BD",x"43",x"1B", -- 0x0500
    x"99",x"4D",x"1D",x"BD",x"4D",x"1B",x"99",x"4E", -- 0x0508
    x"1D",x"BD",x"57",x"1B",x"99",x"4F",x"1D",x"60", -- 0x0510
    x"18",x"29",x"F0",x"4A",x"4A",x"4A",x"4A",x"60", -- 0x0518
    x"A0",x"01",x"A9",x"29",x"99",x"CE",x"1F",x"18", -- 0x0520
    x"69",x"01",x"C8",x"C0",x"06",x"D0",x"F5",x"60", -- 0x0528
    x"98",x"18",x"4A",x"4A",x"4A",x"A8",x"8A",x"18", -- 0x0530
    x"69",x"30",x"99",x"AF",x"1F",x"60",x"A0",x"00", -- 0x0538
    x"A6",x"50",x"F0",x"0B",x"AD",x"BC",x"13",x"99", -- 0x0540
    x"D9",x"1F",x"C8",x"C8",x"CA",x"D0",x"F8",x"C0", -- 0x0548
    x"0A",x"F0",x"0A",x"AD",x"BB",x"13",x"99",x"D9", -- 0x0550
    x"1F",x"C8",x"4C",x"4F",x"15",x"60",x"A5",x"10", -- 0x0558
    x"30",x"12",x"F0",x"10",x"38",x"A5",x"C2",x"C9", -- 0x0560
    x"0C",x"90",x"09",x"A2",x"02",x"B5",x"AA",x"F0", -- 0x0568
    x"04",x"CA",x"10",x"F9",x"60",x"86",x"C1",x"18", -- 0x0570
    x"A5",x"C3",x"69",x"60",x"85",x"C3",x"18",x"4A", -- 0x0578
    x"4A",x"4A",x"4A",x"4A",x"85",x"98",x"A2",x"04", -- 0x0580
    x"86",x"97",x"20",x"54",x"13",x"A4",x"99",x"B9", -- 0x0588
    x"6D",x"00",x"D0",x"04",x"CA",x"10",x"F1",x"60", -- 0x0590
    x"A6",x"C1",x"A9",x"01",x"95",x"AA",x"E6",x"C4", -- 0x0598
    x"A9",x"00",x"85",x"C2",x"95",x"BC",x"A4",x"97", -- 0x05A0
    x"B9",x"68",x"00",x"18",x"69",x"01",x"95",x"B6", -- 0x05A8
    x"0A",x"0A",x"0A",x"95",x"AD",x"A4",x"98",x"B9", -- 0x05B0
    x"60",x"00",x"18",x"69",x"02",x"95",x"B0",x"20", -- 0x05B8
    x"2B",x"12",x"94",x"B3",x"20",x"32",x"12",x"A6", -- 0x05C0
    x"C1",x"95",x"B9",x"20",x"AA",x"16",x"60",x"C6", -- 0x05C8
    x"25",x"D0",x"18",x"A5",x"45",x"85",x"25",x"20", -- 0x05D0
    x"5E",x"15",x"E6",x"C2",x"A9",x"02",x"85",x"C1", -- 0x05D8
    x"AA",x"B5",x"AA",x"D0",x"07",x"C6",x"C1",x"A5", -- 0x05E0
    x"C1",x"10",x"F5",x"60",x"B5",x"BC",x"C9",x"07", -- 0x05E8
    x"D0",x"2D",x"20",x"AA",x"16",x"20",x"9E",x"16", -- 0x05F0
    x"B4",x"B3",x"B1",x"BF",x"38",x"C9",x"2E",x"90", -- 0x05F8
    x"07",x"C9",x"3E",x"B0",x"03",x"4C",x"0F",x"16", -- 0x0600
    x"B4",x"B3",x"AD",x"BB",x"13",x"91",x"BF",x"F6", -- 0x0608
    x"AD",x"B5",x"AD",x"C9",x"A8",x"F0",x"35",x"E6", -- 0x0610
    x"C2",x"20",x"9E",x"16",x"4C",x"29",x"16",x"F6", -- 0x0618
    x"AD",x"E6",x"C2",x"B5",x"AD",x"18",x"4A",x"4A", -- 0x0620
    x"4A",x"95",x"B6",x"B4",x"AD",x"20",x"10",x"12", -- 0x0628
    x"95",x"BC",x"20",x"9E",x"16",x"20",x"C0",x"16", -- 0x0630
    x"20",x"DA",x"16",x"B4",x"B3",x"B1",x"BF",x"4C", -- 0x0638
    x"51",x"16",x"B4",x"B3",x"BD",x"61",x"1B",x"91", -- 0x0640
    x"BF",x"4C",x"E5",x"15",x"A9",x"00",x"95",x"AA", -- 0x0648
    x"60",x"38",x"C9",x"2E",x"90",x"EC",x"C9",x"3E", -- 0x0650
    x"B0",x"E8",x"85",x"56",x"38",x"E9",x"2E",x"85", -- 0x0658
    x"57",x"0A",x"0A",x"0A",x"18",x"75",x"BC",x"85", -- 0x0660
    x"58",x"A8",x"B9",x"70",x"1D",x"B4",x"B9",x"39", -- 0x0668
    x"28",x"14",x"D0",x"09",x"A5",x"56",x"B4",x"B3", -- 0x0670
    x"91",x"BF",x"4C",x"E5",x"15",x"B9",x"2C",x"14", -- 0x0678
    x"85",x"5A",x"A5",x"58",x"A8",x"18",x"69",x"02", -- 0x0680
    x"85",x"5B",x"B9",x"70",x"1D",x"25",x"5A",x"99", -- 0x0688
    x"70",x"1D",x"C8",x"C4",x"5B",x"D0",x"F3",x"A9", -- 0x0690
    x"00",x"95",x"AA",x"4C",x"74",x"16",x"B5",x"AD", -- 0x0698
    x"20",x"00",x"12",x"86",x"BF",x"84",x"C0",x"A6", -- 0x06A0
    x"C1",x"60",x"8A",x"0A",x"0A",x"0A",x"A8",x"18", -- 0x06A8
    x"69",x"08",x"8D",x"BC",x"16",x"A9",x"00",x"99", -- 0x06B0
    x"E8",x"1F",x"C8",x"C0",x"00",x"D0",x"F8",x"60", -- 0x06B8
    x"8A",x"0A",x"0A",x"0A",x"18",x"75",x"BC",x"A8", -- 0x06C0
    x"B5",x"B9",x"AA",x"BD",x"28",x"14",x"99",x"E8", -- 0x06C8
    x"1F",x"88",x"A9",x"00",x"99",x"E8",x"1F",x"A6", -- 0x06D0
    x"C1",x"60",x"B5",x"B6",x"C9",x"14",x"D0",x"17", -- 0x06D8
    x"38",x"B5",x"B0",x"C5",x"00",x"90",x"10",x"A5", -- 0x06E0
    x"00",x"69",x"03",x"D5",x"B0",x"90",x"08",x"A9", -- 0x06E8
    x"00",x"95",x"AA",x"A9",x"80",x"85",x"10",x"A5", -- 0x06F0
    x"11",x"F0",x"25",x"30",x"23",x"B5",x"B0",x"C5", -- 0x06F8
    x"03",x"D0",x"1D",x"B5",x"AD",x"C5",x"04",x"D0", -- 0x0700
    x"17",x"A9",x"00",x"95",x"AA",x"A9",x"80",x"85", -- 0x0708
    x"11",x"20",x"9E",x"16",x"B4",x"B3",x"AD",x"BB", -- 0x0710
    x"13",x"91",x"BF",x"68",x"68",x"4C",x"E5",x"15", -- 0x0718
    x"60",x"20",x"D4",x"17",x"20",x"02",x"18",x"A9", -- 0x0720
    x"F0",x"8D",x"05",x"90",x"85",x"13",x"A2",x"0A", -- 0x0728
    x"BD",x"64",x"1B",x"9D",x"44",x"1E",x"CA",x"10", -- 0x0730
    x"F7",x"A2",x"07",x"BD",x"6F",x"1B",x"9D",x"84", -- 0x0738
    x"1E",x"CA",x"10",x"F7",x"A2",x"10",x"BD",x"77", -- 0x0740
    x"1B",x"9D",x"AA",x"1E",x"CA",x"10",x"F7",x"A2", -- 0x0748
    x"0B",x"BD",x"88",x"1B",x"9D",x"EB",x"1E",x"CA", -- 0x0750
    x"10",x"F7",x"A2",x"04",x"BD",x"94",x"1B",x"9D", -- 0x0758
    x"A9",x"1F",x"CA",x"10",x"F7",x"20",x"B4",x"14", -- 0x0760
    x"A9",x"00",x"8D",x"23",x"02",x"A9",x"18",x"85", -- 0x0768
    x"F0",x"A9",x"80",x"85",x"11",x"AD",x"23",x"02", -- 0x0770
    x"18",x"69",x"30",x"8D",x"F8",x"1E",x"20",x"77", -- 0x0778
    x"1A",x"A5",x"11",x"C9",x"01",x"F0",x"2B",x"A5", -- 0x0780
    x"02",x"F0",x"13",x"EE",x"23",x"02",x"AD",x"23", -- 0x0788
    x"02",x"C9",x"0A",x"D0",x"02",x"A9",x"00",x"8D", -- 0x0790
    x"23",x"02",x"A9",x"18",x"85",x"F0",x"A2",x"FF", -- 0x0798
    x"A0",x"FF",x"88",x"D0",x"FD",x"CA",x"D0",x"F8", -- 0x07A0
    x"C6",x"F0",x"D0",x"C9",x"20",x"0B",x"1A",x"4C", -- 0x07A8
    x"21",x"17",x"20",x"D4",x"17",x"20",x"E3",x"17", -- 0x07B0
    x"20",x"49",x"10",x"20",x"60",x"10",x"A9",x"03", -- 0x07B8
    x"85",x"50",x"A9",x"00",x"8D",x"21",x"02",x"8D", -- 0x07C0
    x"22",x"02",x"20",x"8E",x"14",x"20",x"37",x"19", -- 0x07C8
    x"20",x"DD",x"1A",x"60",x"20",x"DE",x"17",x"20", -- 0x07D0
    x"ED",x"17",x"20",x"3D",x"10",x"60",x"A9",x"00", -- 0x07D8
    x"4C",x"CF",x"1A",x"A9",x"1E",x"20",x"CF",x"1A", -- 0x07E0
    x"A9",x"1F",x"4C",x"CF",x"1A",x"A9",x"01",x"8D", -- 0x07E8
    x"D5",x"1A",x"A9",x"96",x"20",x"CF",x"1A",x"A9", -- 0x07F0
    x"97",x"20",x"CF",x"1A",x"A9",x"00",x"8D",x"D5", -- 0x07F8
    x"1A",x"60",x"A9",x"20",x"8D",x"D5",x"1A",x"A9", -- 0x0800
    x"1E",x"20",x"CF",x"1A",x"A9",x"1F",x"20",x"CF", -- 0x0808
    x"1A",x"A9",x"00",x"8D",x"D5",x"1A",x"60",x"C6", -- 0x0810
    x"27",x"D0",x"5E",x"A5",x"47",x"85",x"27",x"A5", -- 0x0818
    x"10",x"D0",x"19",x"C6",x"50",x"A5",x"50",x"10", -- 0x0820
    x"05",x"68",x"68",x"4C",x"19",x"10",x"20",x"3E", -- 0x0828
    x"15",x"A9",x"00",x"85",x"00",x"85",x"01",x"A9", -- 0x0830
    x"01",x"85",x"10",x"60",x"A2",x"27",x"B5",x"6D", -- 0x0838
    x"F0",x"20",x"8A",x"18",x"4A",x"4A",x"4A",x"A8", -- 0x0840
    x"B9",x"68",x"00",x"C9",x"14",x"D0",x"EC",x"A9", -- 0x0848
    x"00",x"85",x"50",x"A9",x"00",x"85",x"10",x"A2", -- 0x0850
    x"FF",x"20",x"79",x"18",x"CA",x"D0",x"FA",x"4C", -- 0x0858
    x"29",x"18",x"CA",x"10",x"D9",x"A5",x"52",x"C9", -- 0x0860
    x"05",x"F0",x"02",x"E6",x"52",x"20",x"60",x"10", -- 0x0868
    x"20",x"37",x"19",x"20",x"DD",x"1A",x"20",x"49", -- 0x0870
    x"10",x"60",x"C6",x"26",x"D0",x"41",x"A5",x"46", -- 0x0878
    x"85",x"26",x"A5",x"12",x"F0",x"50",x"30",x"38", -- 0x0880
    x"A5",x"0A",x"20",x"2B",x"12",x"AD",x"BB",x"13", -- 0x0888
    x"99",x"00",x"1E",x"C8",x"99",x"00",x"1E",x"A5", -- 0x0890
    x"53",x"D0",x"0B",x"E6",x"0A",x"A5",x"0A",x"C9", -- 0x0898
    x"50",x"F0",x"1D",x"4C",x"AA",x"18",x"C6",x"0A", -- 0x08A0
    x"F0",x"16",x"A5",x"0A",x"20",x"2B",x"12",x"20", -- 0x08A8
    x"32",x"12",x"BD",x"DC",x"13",x"99",x"00",x"1E", -- 0x08B0
    x"C8",x"BD",x"E0",x"13",x"99",x"00",x"1E",x"60", -- 0x08B8
    x"A9",x"00",x"85",x"12",x"85",x"C4",x"A5",x"0A", -- 0x08C0
    x"20",x"2B",x"12",x"AD",x"BB",x"13",x"99",x"00", -- 0x08C8
    x"1E",x"C8",x"99",x"00",x"1E",x"60",x"A5",x"C4", -- 0x08D0
    x"29",x"E0",x"F0",x"E3",x"A9",x"01",x"85",x"12", -- 0x08D8
    x"E6",x"54",x"A6",x"54",x"BD",x"0D",x"11",x"29", -- 0x08E0
    x"07",x"A8",x"B9",x"99",x"1B",x"85",x"55",x"BD", -- 0x08E8
    x"0D",x"11",x"29",x"40",x"85",x"53",x"F0",x"02", -- 0x08F0
    x"A9",x"50",x"85",x"0A",x"60",x"A5",x"12",x"30", -- 0x08F8
    x"23",x"F0",x"21",x"A5",x"0C",x"D0",x"1D",x"38", -- 0x0900
    x"A5",x"03",x"C5",x"0A",x"90",x"16",x"A5",x"0A", -- 0x0908
    x"69",x"03",x"38",x"C5",x"03",x"90",x"0D",x"A9", -- 0x0910
    x"80",x"85",x"12",x"A5",x"55",x"20",x"8E",x"14", -- 0x0918
    x"A9",x"01",x"85",x"C6",x"60",x"A2",x"0F",x"BD", -- 0x0920
    x"70",x"1D",x"9D",x"00",x"02",x"BD",x"B0",x"1D", -- 0x0928
    x"9D",x"10",x"02",x"CA",x"10",x"F1",x"60",x"A2", -- 0x0930
    x"0F",x"BD",x"00",x"02",x"9D",x"70",x"1D",x"9D", -- 0x0938
    x"80",x"1D",x"9D",x"90",x"1D",x"9D",x"A0",x"1D", -- 0x0940
    x"BD",x"10",x"02",x"9D",x"B0",x"1D",x"9D",x"C0", -- 0x0948
    x"1D",x"9D",x"D0",x"1D",x"9D",x"E0",x"1D",x"CA", -- 0x0950
    x"10",x"DF",x"60",x"C6",x"28",x"D0",x"C5",x"A5", -- 0x0958
    x"48",x"85",x"28",x"A5",x"C5",x"F0",x"15",x"C9", -- 0x0960
    x"10",x"D0",x"0D",x"A5",x"C7",x"D0",x"02",x"A9", -- 0x0968
    x"87",x"49",x"08",x"8D",x"0A",x"90",x"85",x"C7", -- 0x0970
    x"C6",x"C5",x"D0",x"05",x"A9",x"00",x"8D",x"0A", -- 0x0978
    x"90",x"A5",x"11",x"F0",x"12",x"30",x"10",x"A5", -- 0x0980
    x"04",x"18",x"69",x"5F",x"38",x"C9",x"C0",x"90", -- 0x0988
    x"06",x"8D",x"0D",x"90",x"4C",x"9C",x"19",x"A9", -- 0x0990
    x"00",x"8D",x"0D",x"90",x"A5",x"C6",x"F0",x"34", -- 0x0998
    x"C9",x"02",x"F0",x"0D",x"C9",x"03",x"F0",x"1F", -- 0x09A0
    x"A9",x"B4",x"8D",x"0C",x"90",x"A9",x"02",x"85", -- 0x09A8
    x"C6",x"EE",x"0C",x"90",x"EE",x"0C",x"90",x"AD", -- 0x09B0
    x"0C",x"90",x"C9",x"E6",x"D0",x"1D",x"A9",x"FA", -- 0x09B8
    x"8D",x"0C",x"90",x"A9",x"03",x"85",x"C6",x"CE", -- 0x09C0
    x"0C",x"90",x"CE",x"0C",x"90",x"AD",x"0C",x"90", -- 0x09C8
    x"C9",x"DC",x"D0",x"07",x"A9",x"00",x"8D",x"0C", -- 0x09D0
    x"90",x"85",x"C6",x"A5",x"12",x"F0",x"21",x"30", -- 0x09D8
    x"1F",x"AD",x"0B",x"90",x"D0",x"0A",x"A9",x"FF", -- 0x09E0
    x"8D",x"0B",x"90",x"A9",x"C8",x"8D",x"0A",x"90", -- 0x09E8
    x"EE",x"0A",x"90",x"CE",x"0B",x"90",x"AD",x"0B", -- 0x09F0
    x"90",x"C9",x"C8",x"F0",x"E9",x"4C",x"05",x"1A", -- 0x09F8
    x"A9",x"00",x"8D",x"0B",x"90",x"A9",x"0F",x"8D", -- 0x0A00
    x"0E",x"90",x"60",x"20",x"B2",x"17",x"A9",x"01", -- 0x0A08
    x"85",x"10",x"85",x"11",x"A9",x"FF",x"85",x"02", -- 0x0A10
    x"A9",x"50",x"85",x"F3",x"4C",x"5A",x"1A",x"20", -- 0x0A18
    x"97",x"10",x"20",x"0D",x"11",x"20",x"3E",x"12", -- 0x0A20
    x"20",x"E6",x"12",x"20",x"CF",x"15",x"20",x"7A", -- 0x0A28
    x"18",x"A5",x"10",x"F0",x"39",x"A5",x"02",x"30", -- 0x0A30
    x"09",x"A5",x"00",x"C9",x"50",x"F0",x"1B",x"4C", -- 0x0A38
    x"46",x"1A",x"A5",x"00",x"F0",x"14",x"C6",x"F3", -- 0x0A40
    x"D0",x"D5",x"A9",x"50",x"85",x"F3",x"A5",x"11", -- 0x0A48
    x"10",x"04",x"A9",x"01",x"85",x"11",x"C6",x"F1", -- 0x0A50
    x"D0",x"C5",x"EE",x"20",x"02",x"AE",x"20",x"02", -- 0x0A58
    x"BD",x"0D",x"11",x"85",x"F1",x"A5",x"02",x"49", -- 0x0A60
    x"FE",x"85",x"02",x"4C",x"1F",x"1A",x"60",x"C6", -- 0x0A68
    x"22",x"D0",x"4A",x"A5",x"42",x"85",x"22",x"A9", -- 0x0A70
    x"00",x"8D",x"20",x"91",x"AD",x"21",x"91",x"AA", -- 0x0A78
    x"A0",x"FF",x"AD",x"11",x"91",x"29",x"10",x"F0", -- 0x0A80
    x"1B",x"A0",x"01",x"A9",x"7F",x"8D",x"22",x"91", -- 0x0A88
    x"AD",x"20",x"91",x"29",x"80",x"F0",x"0D",x"8A", -- 0x0A90
    x"29",x"40",x"F0",x"08",x"A0",x"FF",x"8A",x"29", -- 0x0A98
    x"02",x"F0",x"01",x"C8",x"84",x"02",x"A5",x"11", -- 0x0AA0
    x"30",x"14",x"D0",x"11",x"A0",x"01",x"AD",x"11", -- 0x0AA8
    x"91",x"29",x"20",x"F0",x"06",x"8A",x"29",x"01", -- 0x0AB0
    x"F0",x"01",x"60",x"84",x"11",x"60",x"AD",x"11", -- 0x0AB8
    x"91",x"29",x"20",x"F0",x"F8",x"8A",x"29",x"01", -- 0x0AC0
    x"F0",x"F3",x"A9",x"00",x"85",x"11",x"60",x"8D", -- 0x0AC8
    x"D8",x"1A",x"A0",x"00",x"A9",x"00",x"99",x"00", -- 0x0AD0
    x"00",x"C8",x"D0",x"FA",x"60",x"A2",x"02",x"18", -- 0x0AD8
    x"A9",x"2E",x"9D",x"65",x"1F",x"E8",x"69",x"01", -- 0x0AE0
    x"9D",x"65",x"1F",x"E8",x"E8",x"E8",x"E8",x"69", -- 0x0AE8
    x"01",x"C9",x"36",x"D0",x"ED",x"18",x"A2",x"02", -- 0x0AF0
    x"9D",x"7A",x"1F",x"E8",x"69",x"01",x"9D",x"7A", -- 0x0AF8
    x"1F",x"E8",x"E8",x"E8",x"E8",x"69",x"01",x"C9", -- 0x0B00
    x"3E",x"D0",x"ED",x"60",x"03",x"02",x"02",x"01", -- 0x0B08
    x"01",x"FE",x"18",x"FE",x"FE",x"EC",x"FE",x"FE", -- 0x0B10
    x"FE",x"FE",x"FE",x"FE",x"38",x"FE",x"FE",x"EC", -- 0x0B18
    x"FE",x"E0",x"FE",x"FE",x"FE",x"E6",x"78",x"06", -- 0x0B20
    x"06",x"EC",x"C0",x"E0",x"06",x"E6",x"E6",x"E6", -- 0x0B28
    x"18",x"FE",x"1E",x"FE",x"FE",x"FE",x"0C",x"FE", -- 0x0B30
    x"FE",x"E6",x"18",x"E0",x"1E",x"FE",x"06",x"E6", -- 0x0B38
    x"7E",x"E6",x"FE",x"E6",x"18",x"E0",x"06",x"0C", -- 0x0B40
    x"06",x"E6",x"30",x"E6",x"06",x"FE",x"FE",x"FE", -- 0x0B48
    x"FE",x"0C",x"FE",x"FE",x"60",x"FE",x"06",x"FE", -- 0x0B50
    x"FE",x"FE",x"FE",x"0C",x"FE",x"FE",x"C0",x"FE", -- 0x0B58
    x"06",x"7D",x"7E",x"7F",x"01",x"0C",x"09",x"05", -- 0x0B60
    x"0E",x"20",x"02",x"0C",x"09",x"14",x"1A",x"28", -- 0x0B68
    x"03",x"29",x"20",x"31",x"39",x"38",x"31",x"14", -- 0x0B70
    x"05",x"0E",x"13",x"0F",x"12",x"20",x"14",x"05", -- 0x0B78
    x"03",x"08",x"0E",x"0F",x"0C",x"0F",x"07",x"19", -- 0x0B80
    x"13",x"05",x"0C",x"05",x"03",x"14",x"20",x"0C", -- 0x0B88
    x"05",x"16",x"05",x"0C",x"13",x"03",x"0F",x"12", -- 0x0B90
    x"05",x"05",x"10",x"15",x"20",x"25",x"30",x"40", -- 0x0B98
    x"50",x"FF",x"EA",x"C3",x"9C",x"75",x"4E",x"38", -- 0x0BA0
    x"27",x"10",x"08",x"06",x"06",x"05",x"04",x"03", -- 0x0BA8
    x"02",x"02",x"01",x"00",x"00",x"FF",x"EF",x"EF", -- 0x0BB0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"4D", -- 0x0BB8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0BC0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"49", -- 0x0BC8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0BD0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"4D", -- 0x0BD8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"F7",x"EF",x"EF", -- 0x0BE0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"4D", -- 0x0BE8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0BF0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"49", -- 0x0BF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C00
    x"18",x"3C",x"7E",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C08
    x"06",x"0F",x"1F",x"3F",x"3F",x"3F",x"3F",x"3F", -- 0x0C10
    x"01",x"03",x"07",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x0C18
    x"00",x"00",x"01",x"03",x"03",x"03",x"03",x"03", -- 0x0C20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C28
    x"00",x"00",x"80",x"C0",x"C0",x"C0",x"C0",x"C0", -- 0x0C30
    x"80",x"C0",x"E0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x0C38
    x"60",x"F0",x"F8",x"FC",x"FC",x"FC",x"FC",x"FC", -- 0x0C40
    x"18",x"7E",x"FF",x"99",x"FF",x"24",x"5A",x"81", -- 0x0C48
    x"06",x"1F",x"3F",x"26",x"3F",x"19",x"26",x"10", -- 0x0C50
    x"01",x"07",x"0F",x"09",x"0F",x"02",x"05",x"08", -- 0x0C58
    x"00",x"01",x"03",x"02",x"03",x"01",x"02",x"01", -- 0x0C60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C68
    x"00",x"80",x"C0",x"40",x"C0",x"80",x"40",x"80", -- 0x0C70
    x"80",x"E0",x"F0",x"90",x"F0",x"40",x"A0",x"10", -- 0x0C78
    x"60",x"F8",x"FC",x"64",x"FC",x"98",x"64",x"08", -- 0x0C80
    x"42",x"24",x"3C",x"5A",x"FF",x"BD",x"A5",x"24", -- 0x0C88
    x"10",x"09",x"2F",x"36",x"3F",x"0F",x"10",x"20", -- 0x0C90
    x"04",x"02",x"03",x"05",x"0F",x"0B",x"0A",x"02", -- 0x0C98
    x"01",x"00",x"02",x"03",x"03",x"00",x"01",x"02", -- 0x0CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CA8
    x"80",x"00",x"40",x"C0",x"C0",x"00",x"80",x"40", -- 0x0CB0
    x"20",x"40",x"C0",x"A0",x"F0",x"D0",x"50",x"40", -- 0x0CB8
    x"08",x"90",x"F4",x"6C",x"FC",x"F0",x"08",x"04", -- 0x0CC0
    x"18",x"3C",x"7E",x"DB",x"FF",x"5A",x"81",x"42", -- 0x0CC8
    x"06",x"0F",x"1F",x"36",x"3F",x"0F",x"10",x"20", -- 0x0CD0
    x"01",x"03",x"07",x"0D",x"0F",x"05",x"08",x"04", -- 0x0CD8
    x"00",x"00",x"01",x"03",x"03",x"00",x"01",x"02", -- 0x0CE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CE8
    x"00",x"00",x"80",x"C0",x"C0",x"00",x"80",x"40", -- 0x0CF0
    x"80",x"C0",x"E0",x"B0",x"F0",x"A0",x"10",x"20", -- 0x0CF8
    x"60",x"F0",x"F8",x"6C",x"FC",x"F0",x"08",x"04", -- 0x0D00
    x"00",x"18",x"7E",x"FF",x"7E",x"18",x"24",x"42", -- 0x0D08
    x"06",x"1F",x"3F",x"3F",x"1F",x"06",x"09",x"10", -- 0x0D10
    x"00",x"01",x"07",x"0F",x"07",x"01",x"02",x"04", -- 0x0D18
    x"00",x"01",x"03",x"03",x"01",x"00",x"00",x"01", -- 0x0D20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D28
    x"00",x"80",x"C0",x"C0",x"80",x"00",x"00",x"80", -- 0x0D30
    x"00",x"80",x"E0",x"F0",x"E0",x"80",x"40",x"20", -- 0x0D38
    x"60",x"F8",x"FC",x"FC",x"F8",x"60",x"90",x"08", -- 0x0D40
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0D48
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0D50
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0D58
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0D60
    x"FE",x"FE",x"E6",x"E6",x"E6",x"E6",x"FE",x"FE", -- 0x0D68
    x"03",x"0F",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x0D70
    x"C0",x"F0",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x0D78
    x"03",x"0F",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x0D80
    x"C0",x"F0",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x0D88
    x"03",x"0F",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x0D90
    x"C0",x"F0",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x0D98
    x"03",x"0F",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x0DA0
    x"C0",x"F0",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x0DA8
    x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F8",x"F8", -- 0x0DB0
    x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1F",x"1F", -- 0x0DB8
    x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F8",x"F8", -- 0x0DC0
    x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1F",x"1F", -- 0x0DC8
    x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F8",x"F8", -- 0x0DD0
    x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1F",x"1F", -- 0x0DD8
    x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F8",x"F8", -- 0x0DE0
    x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1F",x"1F", -- 0x0DE8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0DF0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"4D", -- 0x0DF8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E00
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E08
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E10
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E18
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E20
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E28
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E30
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E38
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E40
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E48
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E50
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E58
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E60
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E68
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E70
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E78
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E80
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E88
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E90
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0E98
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0EA0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0EA8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0EB0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0EB8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0EC0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0EC8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0ED0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0ED8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0EE0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0EE8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0EF0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0EF8
    x"A9",x"A0",x"85",x"01",x"A9",x"00",x"85",x"00", -- 0x0F00
    x"85",x"02",x"A9",x"10",x"85",x"03",x"A0",x"00", -- 0x0F08
    x"B1",x"00",x"91",x"02",x"C8",x"D0",x"F9",x"E6", -- 0x0F10
    x"01",x"E6",x"03",x"A5",x"01",x"C9",x"AE",x"D0", -- 0x0F18
    x"EF",x"4C",x"0C",x"10",x"A9",x"60",x"85",x"01", -- 0x0F20
    x"A0",x"00",x"B1",x"00",x"91",x"02",x"C8",x"D0", -- 0x0F28
    x"F9",x"E6",x"01",x"E6",x"03",x"A5",x"01",x"C9", -- 0x0F30
    x"66",x"D0",x"EF",x"60",x"18",x"A2",x"00",x"A0", -- 0x0F38
    x"10",x"20",x"9C",x"FF",x"A9",x"01",x"85",x"2B", -- 0x0F40
    x"A9",x"10",x"85",x"2C",x"60",x"A9",x"00",x"85", -- 0x0F48
    x"2D",x"A9",x"1E",x"85",x"2E",x"60",x"EF",x"EF", -- 0x0F50
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0F58
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0F60
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0F68
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0F70
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0F78
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0F80
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"4D", -- 0x0F88
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0F90
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"4D", -- 0x0F98
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0FA0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"4D", -- 0x0FA8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0FB0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"4D", -- 0x0FB8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0FC0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"4D", -- 0x0FC8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0FD0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"09", -- 0x0FD8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0FE0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"09", -- 0x0FE8
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"EF", -- 0x0FF0
    x"FF",x"FF",x"EF",x"EF",x"FF",x"FF",x"EF",x"49"  -- 0x0FF8
    
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
