-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity cart_rom is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of cart_rom is


  type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"09",x"A0",x"F9",x"BA",x"41",x"30",x"C3",x"C2", -- 0x0000 -- 43 --41
    x"CD",x"D8",x"20",x"8D",x"FD",x"20",x"8A",x"FF", -- 0x0008
    x"20",x"F9",x"FD",x"A9",x"1E",x"8D",x"88",x"02", -- 0x0010
    x"20",x"18",x"E5",x"20",x"5B",x"E4",x"20",x"A4", -- 0x0018
    x"E3",x"78",x"A2",x"FF",x"9A",x"58",x"20",x"7D", -- 0x0020
    x"A1",x"20",x"5A",x"BA",x"20",x"AA",x"A1",x"A9", -- 0x0028
    x"00",x"85",x"F7",x"85",x"F8",x"85",x"F9",x"20", -- 0x0030
    x"B8",x"A1",x"20",x"1B",x"A2",x"20",x"F0",x"A1", -- 0x0038
    x"20",x"C1",x"B4",x"A5",x"42",x"F0",x"08",x"AD", -- 0x0040
    x"0E",x"90",x"09",x"0F",x"8D",x"0E",x"90",x"20", -- 0x0048
    x"1C",x"A4",x"20",x"1C",x"A4",x"20",x"9A",x"A5", -- 0x0050
    x"20",x"61",x"A4",x"A5",x"1E",x"D0",x"08",x"A6", -- 0x0058
    x"20",x"E0",x"02",x"D0",x"0D",x"F0",x"29",x"A5", -- 0x0060
    x"31",x"F0",x"3D",x"A5",x"3E",x"F0",x"E0",x"20", -- 0x0068
    x"F2",x"B4",x"C6",x"3E",x"A5",x"3E",x"C9",x"D0", -- 0x0070
    x"B0",x"D5",x"A6",x"20",x"E0",x"02",x"D0",x"10", -- 0x0078
    x"C9",x"CF",x"D0",x"05",x"AD",x"A6",x"1D",x"85", -- 0x0080
    x"04",x"A5",x"04",x"CD",x"A6",x"1D",x"F0",x"BF", -- 0x0088
    x"A9",x"00",x"85",x"3E",x"85",x"65",x"A5",x"1E", -- 0x0090
    x"F0",x"26",x"A5",x"42",x"D0",x"07",x"A9",x"00", -- 0x0098
    x"85",x"31",x"4C",x"4F",x"A0",x"4C",x"3D",x"A0", -- 0x00A0
    x"A9",x"00",x"85",x"3E",x"78",x"A9",x"68",x"85", -- 0x00A8
    x"35",x"85",x"36",x"A9",x"03",x"85",x"39",x"85", -- 0x00B0
    x"3A",x"58",x"20",x"BB",x"B3",x"4C",x"37",x"A0", -- 0x00B8
    x"A5",x"24",x"C5",x"F9",x"90",x"12",x"D0",x"1C", -- 0x00C0
    x"A5",x"23",x"C5",x"F8",x"90",x"0A",x"D0",x"14", -- 0x00C8
    x"A5",x"22",x"C5",x"F7",x"90",x"02",x"D0",x"0C", -- 0x00D0
    x"A5",x"F7",x"85",x"22",x"A5",x"F8",x"85",x"23", -- 0x00D8
    x"A5",x"F9",x"85",x"24",x"A9",x"00",x"85",x"42", -- 0x00E0
    x"C6",x"1F",x"C6",x"81",x"10",x"02",x"E6",x"81", -- 0x00E8
    x"C6",x"20",x"20",x"94",x"B5",x"A2",x"05",x"86", -- 0x00F0
    x"BE",x"20",x"8E",x"B9",x"C6",x"BE",x"D0",x"F9", -- 0x00F8
    x"4C",x"29",x"A0",x"A4",x"35",x"F0",x"18",x"B9", -- 0x0100
    x"91",x"BE",x"8D",x"0A",x"90",x"D0",x"04",x"85", -- 0x0108
    x"35",x"F0",x"0C",x"C6",x"39",x"D0",x"08",x"C8", -- 0x0110
    x"84",x"35",x"B9",x"20",x"BF",x"85",x"39",x"A4", -- 0x0118
    x"36",x"F0",x"18",x"B9",x"91",x"BE",x"8D",x"0B", -- 0x0120
    x"90",x"D0",x"04",x"85",x"36",x"F0",x"0C",x"C6", -- 0x0128
    x"3A",x"D0",x"08",x"C8",x"84",x"36",x"B9",x"20", -- 0x0130
    x"BF",x"85",x"3A",x"A4",x"37",x"F0",x"18",x"B9", -- 0x0138
    x"91",x"BE",x"8D",x"0C",x"90",x"D0",x"04",x"85", -- 0x0140
    x"37",x"F0",x"0C",x"C6",x"3B",x"D0",x"08",x"C8", -- 0x0148
    x"84",x"37",x"B9",x"20",x"BF",x"85",x"3B",x"A4", -- 0x0150
    x"38",x"F0",x"18",x"B9",x"91",x"BE",x"8D",x"0D", -- 0x0158
    x"90",x"D0",x"04",x"85",x"38",x"F0",x"0C",x"C6", -- 0x0160
    x"3C",x"D0",x"08",x"C8",x"84",x"38",x"B9",x"20", -- 0x0168
    x"BF",x"85",x"3C",x"2C",x"24",x"91",x"68",x"A8", -- 0x0170
    x"68",x"AA",x"68",x"58",x"40",x"A9",x"4C",x"8D", -- 0x0178
    x"5C",x"1D",x"A9",x"00",x"85",x"22",x"85",x"23", -- 0x0180
    x"85",x"24",x"A9",x"80",x"8D",x"91",x"02",x"A2", -- 0x0188
    x"0F",x"BD",x"F8",x"A3",x"9D",x"00",x"90",x"CA", -- 0x0190
    x"10",x"F7",x"20",x"B6",x"A3",x"78",x"A9",x"03", -- 0x0198
    x"8D",x"14",x"03",x"A9",x"A1",x"8D",x"15",x"03", -- 0x01A0
    x"58",x"60",x"A9",x"04",x"85",x"1E",x"A2",x"00", -- 0x01A8
    x"86",x"42",x"86",x"1F",x"E8",x"86",x"81",x"60", -- 0x01B0
    x"A5",x"1F",x"29",x"03",x"85",x"20",x"E6",x"1F", -- 0x01B8
    x"A9",x"10",x"A6",x"20",x"F0",x"05",x"A2",x"0E", -- 0x01C0
    x"0A",x"D0",x"02",x"A2",x"6A",x"8D",x"0E",x"90", -- 0x01C8
    x"8E",x"0F",x"90",x"A9",x"0F",x"85",x"26",x"A2", -- 0x01D0
    x"00",x"86",x"3E",x"86",x"B0",x"86",x"28",x"86", -- 0x01D8
    x"32",x"86",x"3D",x"A2",x"03",x"A9",x"00",x"95", -- 0x01E0
    x"35",x"9D",x"0A",x"90",x"CA",x"10",x"F8",x"60", -- 0x01E8
    x"A2",x"FF",x"8E",x"A4",x"03",x"E8",x"8E",x"5F", -- 0x01F0
    x"1D",x"8E",x"3C",x"03",x"8E",x"56",x"03",x"A9", -- 0x01F8
    x"21",x"8D",x"70",x"03",x"A9",x"9F",x"8D",x"8A", -- 0x0200
    x"03",x"A9",x"FF",x"85",x"2E",x"A9",x"00",x"8D", -- 0x0208
    x"24",x"1D",x"A2",x"05",x"9D",x"44",x"1D",x"CA", -- 0x0210
    x"10",x"FA",x"60",x"A2",x"19",x"A9",x"FF",x"9D", -- 0x0218
    x"3C",x"03",x"9D",x"A4",x"03",x"A9",x"00",x"9D", -- 0x0220
    x"24",x"1D",x"CA",x"D0",x"F0",x"A9",x"64",x"85", -- 0x0228
    x"03",x"A4",x"20",x"F0",x"0C",x"88",x"F0",x"06", -- 0x0230
    x"88",x"D0",x"09",x"4C",x"6A",x"A3",x"4C",x"09", -- 0x0238
    x"A3",x"4C",x"C5",x"A2",x"20",x"AA",x"A3",x"A9", -- 0x0240
    x"7C",x"85",x"03",x"A9",x"36",x"85",x"A3",x"A9", -- 0x0248
    x"31",x"A4",x"1F",x"C0",x"0F",x"90",x"02",x"A9", -- 0x0250
    x"41",x"85",x"A4",x"A9",x"03",x"8D",x"71",x"1D", -- 0x0258
    x"A9",x"00",x"8D",x"6F",x"03",x"85",x"64",x"A0", -- 0x0260
    x"05",x"99",x"74",x"00",x"88",x"10",x"FA",x"A0", -- 0x0268
    x"0A",x"84",x"B3",x"B9",x"BA",x"A2",x"20",x"AD", -- 0x0270
    x"B2",x"20",x"C6",x"B1",x"20",x"AD",x"A2",x"C0", -- 0x0278
    x"06",x"D0",x"F0",x"A9",x"26",x"85",x"A3",x"A5", -- 0x0280
    x"A4",x"E9",x"10",x"85",x"A4",x"85",x"7D",x"B9", -- 0x0288
    x"BA",x"A2",x"20",x"AD",x"B2",x"20",x"BB",x"B1", -- 0x0290
    x"20",x"AD",x"A2",x"10",x"F2",x"A9",x"80",x"85", -- 0x0298
    x"7F",x"A9",x"28",x"85",x"7E",x"A2",x"19",x"86", -- 0x02A0
    x"34",x"E8",x"86",x"31",x"60",x"A5",x"A3",x"18", -- 0x02A8
    x"69",x"04",x"85",x"A3",x"A4",x"B3",x"88",x"84", -- 0x02B0
    x"B3",x"60",x"5A",x"58",x"56",x"54",x"52",x"50", -- 0x02B8
    x"4E",x"5F",x"5E",x"5D",x"5C",x"20",x"AA",x"A3", -- 0x02C0
    x"A2",x"00",x"86",x"60",x"8E",x"89",x"03",x"E8", -- 0x02C8
    x"86",x"64",x"E8",x"86",x"5E",x"E8",x"86",x"62", -- 0x02D0
    x"A2",x"06",x"8E",x"70",x"1D",x"8E",x"71",x"1D", -- 0x02D8
    x"A2",x"18",x"86",x"63",x"86",x"31",x"86",x"61", -- 0x02E0
    x"E8",x"86",x"34",x"A9",x"00",x"A0",x"05",x"84", -- 0x02E8
    x"65",x"99",x"74",x"00",x"88",x"10",x"FA",x"A9", -- 0x02F0
    x"07",x"A0",x"59",x"99",x"24",x"96",x"88",x"10", -- 0x02F8
    x"FA",x"A9",x"84",x"85",x"03",x"20",x"52",x"B0", -- 0x0300
    x"60",x"A0",x"B0",x"8C",x"F0",x"03",x"A0",x"01", -- 0x0308
    x"8C",x"71",x"1D",x"A0",x"03",x"A5",x"1F",x"C9", -- 0x0310
    x"09",x"90",x"06",x"C8",x"C9",x"11",x"90",x"01", -- 0x0318
    x"C8",x"84",x"66",x"A0",x"0A",x"84",x"34",x"84", -- 0x0320
    x"31",x"8C",x"70",x"1D",x"B9",x"5F",x"A3",x"99", -- 0x0328
    x"56",x"03",x"A9",x"00",x"99",x"3C",x"03",x"88", -- 0x0330
    x"D0",x"F2",x"C8",x"B9",x"5E",x"A3",x"99",x"71", -- 0x0338
    x"03",x"A9",x"40",x"99",x"8B",x"03",x"A9",x"00", -- 0x0340
    x"99",x"7D",x"03",x"A9",x"FF",x"99",x"6E",x"1D", -- 0x0348
    x"88",x"10",x"E8",x"98",x"A0",x"07",x"99",x"66", -- 0x0350
    x"1D",x"88",x"10",x"FA",x"30",x"4C",x"10",x"34", -- 0x0358
    x"08",x"08",x"10",x"0C",x"0C",x"0C",x"10",x"0C", -- 0x0360
    x"0C",x"0C",x"A9",x"02",x"85",x"34",x"A2",x"FF", -- 0x0368
    x"8E",x"3D",x"03",x"8E",x"72",x"03",x"E8",x"8E", -- 0x0370
    x"A1",x"1D",x"8E",x"A2",x"1D",x"A9",x"41",x"8D", -- 0x0378
    x"57",x"03",x"A9",x"04",x"8D",x"A9",x"1D",x"A9", -- 0x0380
    x"20",x"8D",x"AA",x"1D",x"A9",x"24",x"85",x"5E", -- 0x0388
    x"A9",x"58",x"85",x"5F",x"A9",x"0C",x"A6",x"1F", -- 0x0390
    x"E0",x"03",x"F0",x"02",x"A9",x"10",x"8D",x"A6", -- 0x0398
    x"1D",x"A9",x"11",x"85",x"31",x"A9",x"02",x"8D", -- 0x03A0
    x"2E",x"1D",x"20",x"DF",x"A3",x"20",x"08",x"A4", -- 0x03A8
    x"20",x"C1",x"B4",x"20",x"F2",x"B4",x"A9",x"11", -- 0x03B0
    x"85",x"A5",x"85",x"A7",x"A9",x"1E",x"85",x"A6", -- 0x03B8
    x"A9",x"96",x"85",x"A8",x"A2",x"C5",x"A0",x"B4", -- 0x03C0
    x"8A",x"91",x"A5",x"A5",x"26",x"91",x"A7",x"CA", -- 0x03C8
    x"98",x"38",x"E9",x"12",x"A8",x"B0",x"F1",x"C6", -- 0x03D0
    x"A5",x"C6",x"A7",x"E0",x"FF",x"D0",x"E7",x"A9", -- 0x03D8
    x"00",x"85",x"A5",x"A9",x"10",x"85",x"A6",x"A9", -- 0x03E0
    x"00",x"A8",x"91",x"A5",x"C8",x"D0",x"FB",x"E6", -- 0x03E8
    x"A6",x"A6",x"A6",x"E0",x"1D",x"D0",x"F3",x"60", -- 0x03F0
    x"09",x"1B",x"92",x"17",x"00",x"FC",x"00",x"00", -- 0x03F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08", -- 0x0400
    x"A9",x"00",x"85",x"A7",x"A9",x"96",x"85",x"A8", -- 0x0408
    x"A0",x"C7",x"A5",x"26",x"91",x"A7",x"88",x"C0", -- 0x0410
    x"FF",x"D0",x"F9",x"60",x"A6",x"42",x"D0",x"03", -- 0x0418
    x"4C",x"6E",x"BA",x"AD",x"56",x"03",x"D0",x"38", -- 0x0420
    x"20",x"D8",x"B0",x"24",x"B0",x"10",x"03",x"20", -- 0x0428
    x"52",x"B6",x"18",x"A5",x"B1",x"6D",x"70",x"03", -- 0x0430
    x"C9",x"01",x"B0",x"04",x"A9",x"01",x"D0",x"06", -- 0x0438
    x"C9",x"40",x"90",x"02",x"A9",x"40",x"8D",x"70", -- 0x0440
    x"03",x"18",x"A5",x"B2",x"6D",x"8A",x"03",x"C5", -- 0x0448
    x"03",x"B0",x"04",x"A5",x"03",x"D0",x"06",x"C9", -- 0x0450
    x"A0",x"90",x"02",x"A9",x"A0",x"8D",x"8A",x"03", -- 0x0458
    x"60",x"20",x"93",x"B6",x"A9",x"05",x"85",x"B4", -- 0x0460
    x"A6",x"B4",x"BD",x"44",x"1D",x"F0",x"33",x"BD", -- 0x0468
    x"4A",x"1D",x"85",x"A3",x"BD",x"50",x"1D",x"85", -- 0x0470
    x"A4",x"20",x"4C",x"A5",x"98",x"30",x"23",x"A6", -- 0x0478
    x"B4",x"D0",x"05",x"98",x"F0",x"1C",x"D0",x"03", -- 0x0480
    x"98",x"D0",x"17",x"20",x"A1",x"B8",x"A6",x"B4", -- 0x0488
    x"20",x"45",x"B7",x"A9",x"43",x"20",x"AD",x"B2", -- 0x0490
    x"20",x"50",x"B2",x"A6",x"B4",x"A9",x"00",x"9D", -- 0x0498
    x"44",x"1D",x"C6",x"B4",x"10",x"C2",x"A5",x"34", -- 0x04A0
    x"85",x"B4",x"A4",x"B4",x"B9",x"3C",x"03",x"C9", -- 0x04A8
    x"FF",x"F0",x"23",x"B9",x"56",x"03",x"C9",x"44", -- 0x04B0
    x"90",x"06",x"20",x"A1",x"B8",x"4C",x"C3",x"A4", -- 0x04B8
    x"20",x"13",x"B2",x"A4",x"B4",x"20",x"89",x"B1", -- 0x04C0
    x"A4",x"B4",x"B9",x"70",x"03",x"99",x"A4",x"03", -- 0x04C8
    x"B9",x"8A",x"03",x"99",x"BE",x"03",x"C6",x"B4", -- 0x04D0
    x"10",x"D0",x"AD",x"56",x"03",x"D0",x"1A",x"AD", -- 0x04D8
    x"70",x"03",x"85",x"A3",x"AD",x"8A",x"03",x"85", -- 0x04E0
    x"A4",x"20",x"FA",x"A4",x"98",x"30",x"0A",x"F0", -- 0x04E8
    x"08",x"20",x"A1",x"B8",x"A0",x"00",x"20",x"A1", -- 0x04F0
    x"B8",x"60",x"A4",x"34",x"B9",x"3C",x"03",x"30", -- 0x04F8
    x"47",x"BE",x"56",x"03",x"E0",x"35",x"F0",x"40", -- 0x0500
    x"A9",x"04",x"E0",x"38",x"B0",x"01",x"0A",x"85", -- 0x0508
    x"01",x"0A",x"85",x"02",x"B9",x"70",x"03",x"C5", -- 0x0510
    x"A3",x"B0",x"09",x"18",x"65",x"01",x"C5",x"A3", -- 0x0518
    x"B0",x"0C",x"90",x"24",x"A5",x"A3",x"18",x"65", -- 0x0520
    x"01",x"D9",x"70",x"03",x"90",x"1A",x"B9",x"8A", -- 0x0528
    x"03",x"C5",x"A4",x"B0",x"09",x"18",x"65",x"02", -- 0x0530
    x"C5",x"A4",x"B0",x"0F",x"90",x"0A",x"A5",x"A4", -- 0x0538
    x"18",x"65",x"02",x"D9",x"8A",x"03",x"B0",x"03", -- 0x0540
    x"88",x"10",x"B1",x"60",x"A4",x"34",x"B9",x"3C", -- 0x0548
    x"03",x"30",x"43",x"BE",x"56",x"03",x"E0",x"44", -- 0x0550
    x"B0",x"3C",x"E0",x"42",x"F0",x"38",x"E0",x"14", -- 0x0558
    x"F0",x"34",x"E0",x"18",x"F0",x"30",x"E0",x"35", -- 0x0560
    x"F0",x"2C",x"A9",x"04",x"E0",x"38",x"B0",x"01", -- 0x0568
    x"0A",x"85",x"01",x"0A",x"85",x"02",x"B9",x"70", -- 0x0570
    x"03",x"C5",x"A3",x"F0",x"09",x"B0",x"17",x"18", -- 0x0578
    x"65",x"01",x"C5",x"A3",x"90",x"10",x"B9",x"8A", -- 0x0580
    x"03",x"C5",x"A4",x"F0",x"0C",x"B0",x"07",x"18", -- 0x0588
    x"65",x"02",x"C5",x"A4",x"B0",x"03",x"88",x"10", -- 0x0590
    x"B5",x"60",x"A5",x"20",x"29",x"03",x"A8",x"F0", -- 0x0598
    x"09",x"88",x"F0",x"09",x"88",x"F0",x"09",x"4C", -- 0x05A0
    x"E7",x"AE",x"4C",x"D1",x"A5",x"4C",x"00",x"A8", -- 0x05A8
    x"4C",x"D6",x"AA",x"02",x"08",x"0E",x"14",x"1A", -- 0x05B0
    x"20",x"26",x"2C",x"2C",x"26",x"20",x"1A",x"14", -- 0x05B8
    x"0E",x"08",x"02",x"02",x"08",x"0E",x"14",x"1A", -- 0x05C0
    x"20",x"26",x"2C",x"30",x"3C",x"48",x"39",x"3A", -- 0x05C8
    x"3B",x"20",x"52",x"B0",x"A5",x"61",x"F0",x"58", -- 0x05D0
    x"20",x"F5",x"A6",x"AD",x"89",x"03",x"C9",x"30", -- 0x05D8
    x"B0",x"47",x"A5",x"65",x"D0",x"47",x"78",x"A9", -- 0x05E0
    x"77",x"85",x"36",x"A9",x"04",x"85",x"3A",x"58", -- 0x05E8
    x"A9",x"04",x"85",x"65",x"A6",x"62",x"A4",x"63", -- 0x05F0
    x"B9",x"B2",x"A5",x"99",x"70",x"03",x"A5",x"1F", -- 0x05F8
    x"0A",x"C9",x"28",x"90",x"02",x"A9",x"28",x"7D", -- 0x0600
    x"CA",x"A5",x"99",x"8A",x"03",x"BD",x"CD",x"A5", -- 0x0608
    x"99",x"56",x"03",x"A9",x"00",x"99",x"3C",x"03", -- 0x0610
    x"A4",x"63",x"88",x"F0",x"0D",x"C0",x"10",x"F0", -- 0x0618
    x"04",x"C0",x"08",x"D0",x"02",x"C6",x"62",x"84", -- 0x0620
    x"63",x"60",x"84",x"61",x"60",x"C6",x"65",x"60", -- 0x0628
    x"AD",x"14",x"91",x"CD",x"71",x"1D",x"90",x"04", -- 0x0630
    x"A5",x"64",x"F0",x"03",x"20",x"F5",x"A6",x"AD", -- 0x0638
    x"56",x"03",x"F0",x"03",x"4C",x"F2",x"A6",x"A5", -- 0x0640
    x"65",x"F0",x"03",x"4C",x"F2",x"A6",x"78",x"A9", -- 0x0648
    x"01",x"85",x"35",x"A9",x"02",x"85",x"39",x"58", -- 0x0650
    x"A2",x"05",x"A5",x"31",x"C9",x"02",x"F0",x"04", -- 0x0658
    x"C9",x"01",x"D0",x"01",x"AA",x"86",x"65",x"A5", -- 0x0660
    x"5E",x"C9",x"44",x"D0",x"04",x"A9",x"FE",x"D0", -- 0x0668
    x"02",x"A9",x"02",x"85",x"5F",x"A0",x"18",x"B9", -- 0x0670
    x"3C",x"03",x"30",x"4B",x"B9",x"56",x"03",x"C9", -- 0x0678
    x"44",x"B0",x"44",x"84",x"BF",x"20",x"13",x"B2", -- 0x0680
    x"A4",x"BF",x"B9",x"56",x"03",x"49",x"07",x"99", -- 0x0688
    x"56",x"03",x"B9",x"70",x"03",x"18",x"65",x"5F", -- 0x0690
    x"99",x"70",x"03",x"AE",x"14",x"91",x"EC",x"70", -- 0x0698
    x"1D",x"90",x"0E",x"E9",x"03",x"CD",x"70",x"03", -- 0x06A0
    x"B0",x"0E",x"69",x"06",x"CD",x"70",x"03",x"90", -- 0x06A8
    x"07",x"84",x"2F",x"20",x"55",x"B7",x"A4",x"2F", -- 0x06B0
    x"B9",x"70",x"03",x"F0",x"04",x"C9",x"44",x"D0", -- 0x06B8
    x"06",x"85",x"5E",x"A9",x"FF",x"85",x"60",x"88", -- 0x06C0
    x"D0",x"AD",x"A5",x"60",x"F0",x"23",x"A0",x"18", -- 0x06C8
    x"B9",x"56",x"03",x"C9",x"44",x"B0",x"15",x"B9", -- 0x06D0
    x"8A",x"03",x"69",x"06",x"C9",x"A8",x"90",x"09", -- 0x06D8
    x"AD",x"70",x"03",x"99",x"70",x"03",x"AD",x"8A", -- 0x06E0
    x"03",x"99",x"8A",x"03",x"88",x"D0",x"E1",x"84", -- 0x06E8
    x"60",x"60",x"C6",x"65",x"60",x"AD",x"6F",x"03", -- 0x06F0
    x"C9",x"46",x"90",x"01",x"60",x"A5",x"64",x"30", -- 0x06F8
    x"61",x"09",x"80",x"85",x"64",x"A9",x"00",x"8D", -- 0x0700
    x"55",x"03",x"A9",x"3E",x"8D",x"89",x"03",x"A9", -- 0x0708
    x"08",x"8D",x"A3",x"03",x"A9",x"FF",x"85",x"04", -- 0x0710
    x"A2",x"02",x"86",x"05",x"A2",x"20",x"86",x"06", -- 0x0718
    x"A5",x"64",x"C9",x"81",x"F0",x"31",x"AD",x"14", -- 0x0720
    x"91",x"29",x"01",x"F0",x"05",x"85",x"04",x"8D", -- 0x0728
    x"89",x"03",x"AD",x"14",x"91",x"C9",x"A9",x"B0", -- 0x0730
    x"06",x"A9",x"82",x"85",x"64",x"D0",x"18",x"A9", -- 0x0738
    x"00",x"85",x"05",x"A5",x"04",x"0A",x"85",x"04", -- 0x0740
    x"EE",x"A3",x"03",x"A2",x"83",x"AD",x"15",x"91", -- 0x0748
    x"29",x"01",x"F0",x"01",x"E8",x"86",x"64",x"A5", -- 0x0750
    x"64",x"29",x"07",x"AA",x"BD",x"FB",x"A7",x"8D", -- 0x0758
    x"6F",x"03",x"A5",x"04",x"F0",x"54",x"18",x"6D", -- 0x0760
    x"89",x"03",x"8D",x"89",x"03",x"AD",x"A3",x"03", -- 0x0768
    x"18",x"65",x"05",x"8D",x"A3",x"03",x"C9",x"08", -- 0x0770
    x"F0",x"04",x"C9",x"10",x"D0",x"06",x"A5",x"05", -- 0x0778
    x"49",x"FC",x"85",x"05",x"A5",x"64",x"C9",x"84", -- 0x0780
    x"F0",x"10",x"C9",x"81",x"F0",x"42",x"AD",x"89", -- 0x0788
    x"03",x"C9",x"60",x"90",x"04",x"C9",x"F0",x"90", -- 0x0790
    x"5A",x"60",x"AD",x"A3",x"03",x"C9",x"09",x"D0", -- 0x0798
    x"ED",x"AD",x"89",x"03",x"C9",x"30",x"90",x"06", -- 0x07A0
    x"A6",x"04",x"30",x"E2",x"10",x"08",x"C9",x"18", -- 0x07A8
    x"D0",x"DC",x"A6",x"04",x"10",x"D8",x"A9",x"00", -- 0x07B0
    x"85",x"04",x"C6",x"06",x"D0",x"D0",x"EE",x"A3", -- 0x07B8
    x"03",x"A2",x"02",x"AD",x"89",x"03",x"C9",x"30", -- 0x07C0
    x"90",x"02",x"A2",x"FE",x"86",x"04",x"D0",x"BE", -- 0x07C8
    x"AD",x"89",x"03",x"C9",x"03",x"D0",x"04",x"A5", -- 0x07D0
    x"04",x"30",x"0E",x"C9",x"28",x"D0",x"AF",x"A5", -- 0x07D8
    x"04",x"30",x"AB",x"A9",x"82",x"85",x"64",x"A5", -- 0x07E0
    x"04",x"49",x"FE",x"85",x"04",x"A9",x"02",x"85", -- 0x07E8
    x"05",x"D0",x"9B",x"A9",x"00",x"85",x"04",x"85", -- 0x07F0
    x"05",x"85",x"64",x"60",x"04",x"04",x"2C",x"2F", -- 0x07F8
    x"A2",x"01",x"AD",x"56",x"03",x"D0",x"30",x"BD", -- 0x0800
    x"6E",x"1D",x"D0",x"2B",x"BD",x"7D",x"03",x"D0", -- 0x0808
    x"2C",x"AD",x"14",x"91",x"CD",x"F0",x"03",x"90", -- 0x0810
    x"24",x"BD",x"57",x"03",x"C9",x"44",x"B0",x"1D", -- 0x0818
    x"20",x"3D",x"AA",x"BD",x"57",x"03",x"C9",x"08", -- 0x0820
    x"D0",x"13",x"AD",x"14",x"91",x"CD",x"70",x"1D", -- 0x0828
    x"90",x"05",x"A9",x"FF",x"9D",x"6E",x"1D",x"20", -- 0x0830
    x"53",x"A9",x"4C",x"45",x"A8",x"BD",x"7D",x"03", -- 0x0838
    x"F0",x"03",x"20",x"3D",x"AA",x"CA",x"10",x"BA", -- 0x0840
    x"A2",x"01",x"A0",x"07",x"B9",x"59",x"03",x"D9", -- 0x0848
    x"62",x"A3",x"F0",x"0A",x"A9",x"FF",x"85",x"BE", -- 0x0850
    x"C6",x"BE",x"F0",x"48",x"D0",x"FA",x"B9",x"66", -- 0x0858
    x"1D",x"10",x"32",x"AD",x"56",x"03",x"D0",x"16", -- 0x0860
    x"BD",x"57",x"03",x"C9",x"08",x"D0",x"08",x"AD", -- 0x0868
    x"14",x"91",x"CD",x"71",x"1D",x"B0",x"07",x"A9", -- 0x0870
    x"01",x"99",x"66",x"1D",x"90",x"1F",x"BD",x"8B", -- 0x0878
    x"03",x"18",x"79",x"B7",x"A8",x"99",x"8D",x"03", -- 0x0880
    x"BD",x"71",x"03",x"18",x"79",x"AF",x"A8",x"99", -- 0x0888
    x"73",x"03",x"4C",x"A4",x"A8",x"D0",x"06",x"20", -- 0x0890
    x"40",x"A9",x"4C",x"A4",x"A8",x"86",x"BE",x"20", -- 0x0898
    x"BF",x"A8",x"A6",x"BE",x"88",x"10",x"01",x"60", -- 0x08A0
    x"C0",x"03",x"D0",x"A0",x"CA",x"10",x"9D",x"00", -- 0x08A8
    x"F8",x"00",x"08",x"00",x"F8",x"00",x"08",x"E0", -- 0x08B0
    x"F2",x"F2",x"F2",x"E0",x"F2",x"F2",x"F2",x"78", -- 0x08B8
    x"AD",x"0B",x"90",x"30",x"08",x"A9",x"40",x"85", -- 0x08C0
    x"36",x"A9",x"02",x"85",x"3A",x"58",x"18",x"B9", -- 0x08C8
    x"8D",x"03",x"65",x"66",x"C9",x"A0",x"99",x"8D", -- 0x08D0
    x"03",x"90",x"19",x"A9",x"00",x"99",x"66",x"1D", -- 0x08D8
    x"A9",x"10",x"99",x"8D",x"03",x"BD",x"71",x"03", -- 0x08E0
    x"99",x"73",x"03",x"BD",x"8B",x"03",x"38",x"E9", -- 0x08E8
    x"20",x"95",x"5E",x"60",x"C9",x"80",x"B0",x"25", -- 0x08F0
    x"A2",x"00",x"38",x"B9",x"73",x"03",x"ED",x"70", -- 0x08F8
    x"03",x"F0",x"0B",x"10",x"08",x"49",x"FF",x"18", -- 0x0900
    x"69",x"01",x"E8",x"D0",x"01",x"CA",x"86",x"5A", -- 0x0908
    x"A2",x"06",x"DD",x"39",x"A9",x"90",x"03",x"CA", -- 0x0910
    x"D0",x"F8",x"E8",x"86",x"5B",x"A6",x"5C",x"D0", -- 0x0918
    x"14",x"A6",x"5A",x"F0",x"0E",x"30",x"07",x"98", -- 0x0920
    x"AA",x"FE",x"73",x"03",x"D0",x"05",x"98",x"AA", -- 0x0928
    x"DE",x"73",x"03",x"A6",x"5B",x"CA",x"86",x"5C", -- 0x0930
    x"60",x"3C",x"1E",x"14",x"0F",x"0A",x"05",x"00", -- 0x0938
    x"18",x"B9",x"8D",x"03",x"65",x"66",x"99",x"8D", -- 0x0940
    x"03",x"D5",x"5E",x"90",x"05",x"A9",x"FF",x"99", -- 0x0948
    x"66",x"1D",x"60",x"BD",x"6E",x"1D",x"F0",x"55", -- 0x0950
    x"B5",x"67",x"85",x"6B",x"B5",x"69",x"85",x"6C", -- 0x0958
    x"18",x"BD",x"71",x"03",x"69",x"03",x"85",x"6D", -- 0x0960
    x"BD",x"6E",x"1D",x"10",x"41",x"78",x"A9",x"68", -- 0x0968
    x"85",x"36",x"85",x"35",x"A9",x"03",x"85",x"3A", -- 0x0970
    x"85",x"39",x"58",x"A5",x"6D",x"29",x"03",x"A8", -- 0x0978
    x"B9",x"A9",x"B2",x"95",x"07",x"A5",x"6D",x"4A", -- 0x0980
    x"29",x"FE",x"A8",x"18",x"B9",x"5F",x"B1",x"69", -- 0x0988
    x"0E",x"7D",x"8B",x"03",x"95",x"67",x"B9",x"60", -- 0x0990
    x"B1",x"69",x"00",x"95",x"69",x"A9",x"A0",x"FD", -- 0x0998
    x"8B",x"03",x"95",x"0B",x"A9",x"00",x"95",x"09", -- 0x09A0
    x"A9",x"02",x"9D",x"6E",x"1D",x"60",x"C9",x"01", -- 0x09A8
    x"D0",x"33",x"B5",x"09",x"85",x"6E",x"A0",x"00", -- 0x09B0
    x"B5",x"07",x"49",x"FF",x"31",x"6B",x"91",x"6B", -- 0x09B8
    x"C8",x"C4",x"6E",x"D0",x"F3",x"A5",x"6E",x"D5", -- 0x09C0
    x"0B",x"90",x"0D",x"A9",x"00",x"9D",x"6E",x"1D", -- 0x09C8
    x"86",x"BE",x"20",x"DB",x"B4",x"A6",x"BE",x"60", -- 0x09D0
    x"B5",x"0B",x"85",x"6E",x"B5",x"09",x"18",x"69", -- 0x09D8
    x"07",x"95",x"09",x"D0",x"17",x"18",x"B5",x"09", -- 0x09E0
    x"69",x"07",x"D5",x"0B",x"90",x"08",x"A9",x"01", -- 0x09E8
    x"9D",x"6E",x"1D",x"95",x"09",x"60",x"85",x"6E", -- 0x09F0
    x"95",x"09",x"A0",x"00",x"AD",x"56",x"03",x"D0", -- 0x09F8
    x"30",x"AD",x"70",x"03",x"C5",x"6D",x"F0",x"08", -- 0x0A00
    x"B0",x"27",x"69",x"07",x"C5",x"6D",x"90",x"21", -- 0x0A08
    x"84",x"AD",x"AD",x"8A",x"03",x"FD",x"8B",x"03", -- 0x0A10
    x"E9",x"10",x"C5",x"6E",x"F0",x"02",x"B0",x"11", -- 0x0A18
    x"18",x"69",x"0F",x"C5",x"AD",x"90",x"0A",x"86", -- 0x0A20
    x"BE",x"A0",x"00",x"20",x"A1",x"B8",x"A6",x"BE", -- 0x0A28
    x"60",x"B5",x"07",x"11",x"6B",x"91",x"6B",x"C8", -- 0x0A30
    x"C4",x"6E",x"D0",x"F5",x"60",x"BD",x"7D",x"03", -- 0x0A38
    x"D0",x"52",x"AD",x"14",x"91",x"29",x"07",x"E0", -- 0x0A40
    x"01",x"D0",x"03",x"18",x"69",x"07",x"A8",x"B9", -- 0x0A48
    x"C7",x"AA",x"6D",x"70",x"03",x"C9",x"0A",x"10", -- 0x0A50
    x"04",x"A9",x"0A",x"D0",x"06",x"C9",x"2F",x"90", -- 0x0A58
    x"02",x"A9",x"2F",x"9D",x"7B",x"03",x"AD",x"7B", -- 0x0A60
    x"03",x"38",x"ED",x"7C",x"03",x"B0",x"04",x"49", -- 0x0A68
    x"FF",x"69",x"01",x"C9",x"04",x"B0",x"05",x"A9", -- 0x0A70
    x"27",x"9D",x"7B",x"03",x"AD",x"14",x"91",x"29", -- 0x0A78
    x"3F",x"18",x"69",x"30",x"9D",x"95",x"03",x"69", -- 0x0A80
    x"04",x"9D",x"99",x"03",x"BD",x"7B",x"03",x"69", -- 0x0A88
    x"04",x"9D",x"7F",x"03",x"A0",x"00",x"BD",x"71", -- 0x0A90
    x"03",x"DD",x"7B",x"03",x"B0",x"03",x"C8",x"69", -- 0x0A98
    x"03",x"DD",x"7F",x"03",x"90",x"03",x"C8",x"E9", -- 0x0AA0
    x"03",x"9D",x"71",x"03",x"BD",x"8B",x"03",x"DD", -- 0x0AA8
    x"95",x"03",x"B0",x"03",x"C8",x"69",x"03",x"DD", -- 0x0AB0
    x"99",x"03",x"90",x"03",x"C8",x"E9",x"03",x"9D", -- 0x0AB8
    x"8B",x"03",x"98",x"9D",x"7D",x"03",x"60",x"E4", -- 0x0AC0
    x"E4",x"E8",x"EC",x"F0",x"F4",x"F8",x"FC",x"00", -- 0x0AC8
    x"04",x"08",x"0C",x"10",x"14",x"14",x"AE",x"A6", -- 0x0AD0
    x"1D",x"E8",x"8E",x"A7",x"1D",x"BD",x"3E",x"AE", -- 0x0AD8
    x"85",x"A3",x"BD",x"4F",x"AE",x"85",x"A4",x"A9", -- 0x0AE0
    x"71",x"20",x"AD",x"B2",x"20",x"0D",x"B2",x"CE", -- 0x0AE8
    x"A7",x"1D",x"AE",x"A7",x"1D",x"BD",x"3E",x"AE", -- 0x0AF0
    x"85",x"A3",x"BD",x"4F",x"AE",x"85",x"A4",x"A9", -- 0x0AF8
    x"71",x"20",x"AD",x"B2",x"20",x"C6",x"B1",x"AE", -- 0x0B00
    x"A7",x"1D",x"D0",x"E3",x"CE",x"2E",x"1D",x"F0", -- 0x0B08
    x"03",x"4C",x"3D",x"AC",x"A2",x"02",x"A5",x"1F", -- 0x0B10
    x"C9",x"0A",x"90",x"01",x"CA",x"8E",x"2E",x"1D", -- 0x0B18
    x"AD",x"3D",x"03",x"F0",x"08",x"A9",x"00",x"8D", -- 0x0B20
    x"3D",x"03",x"8D",x"A0",x"1D",x"AD",x"57",x"03", -- 0x0B28
    x"C9",x"44",x"90",x"03",x"4C",x"2A",x"AC",x"AD", -- 0x0B30
    x"A0",x"1D",x"F0",x"11",x"C9",x"1C",x"F0",x"04", -- 0x0B38
    x"C9",x"38",x"D0",x"47",x"EE",x"A5",x"1D",x"20", -- 0x0B40
    x"37",x"AC",x"4C",x"8B",x"AB",x"8D",x"A5",x"1D", -- 0x0B48
    x"CE",x"A6",x"1D",x"10",x"05",x"A9",x"00",x"85", -- 0x0B50
    x"31",x"60",x"AD",x"14",x"91",x"29",x"03",x"F0", -- 0x0B58
    x"F9",x"AA",x"BD",x"3A",x"AE",x"8D",x"A8",x"1D", -- 0x0B60
    x"AD",x"14",x"91",x"29",x"01",x"F0",x"02",x"A9", -- 0x0B68
    x"3F",x"8D",x"A1",x"1D",x"AD",x"15",x"91",x"29", -- 0x0B70
    x"01",x"F0",x"02",x"A9",x"7F",x"8D",x"A2",x"1D", -- 0x0B78
    x"AD",x"18",x"91",x"0D",x"19",x"91",x"29",x"01", -- 0x0B80
    x"8D",x"A3",x"1D",x"AE",x"A0",x"1D",x"E0",x"54", -- 0x0B88
    x"90",x"10",x"A9",x"00",x"8D",x"A0",x"1D",x"20", -- 0x0B90
    x"37",x"AC",x"A9",x"C0",x"8D",x"71",x"03",x"4C", -- 0x0B98
    x"2A",x"AC",x"BD",x"E7",x"AD",x"0A",x"4D",x"A1", -- 0x0BA0
    x"1D",x"8D",x"71",x"03",x"E8",x"BD",x"E7",x"AD", -- 0x0BA8
    x"0A",x"0A",x"4D",x"A2",x"1D",x"8D",x"8B",x"03", -- 0x0BB0
    x"E8",x"8E",x"A0",x"1D",x"AD",x"A3",x"1D",x"D0", -- 0x0BB8
    x"14",x"AD",x"71",x"03",x"0A",x"8D",x"A4",x"1D", -- 0x0BC0
    x"AD",x"8B",x"03",x"4A",x"8D",x"71",x"03",x"AD", -- 0x0BC8
    x"A4",x"1D",x"8D",x"8B",x"03",x"AD",x"8B",x"03", -- 0x0BD0
    x"18",x"69",x"18",x"8D",x"8B",x"03",x"AD",x"71", -- 0x0BD8
    x"03",x"18",x"69",x"04",x"8D",x"71",x"03",x"AD", -- 0x0BE0
    x"A8",x"1D",x"18",x"6D",x"A5",x"1D",x"AA",x"BD", -- 0x0BE8
    x"DE",x"AD",x"8D",x"57",x"03",x"AD",x"56",x"03", -- 0x0BF0
    x"D0",x"30",x"A0",x"02",x"B9",x"3C",x"03",x"F0", -- 0x0BF8
    x"29",x"AD",x"71",x"03",x"99",x"70",x"03",x"AD", -- 0x0C00
    x"8B",x"03",x"18",x"69",x"11",x"99",x"8A",x"03", -- 0x0C08
    x"A9",x"42",x"99",x"56",x"03",x"20",x"60",x"AE", -- 0x0C10
    x"78",x"A9",x"75",x"85",x"36",x"A9",x"28",x"85", -- 0x0C18
    x"3A",x"A9",x"51",x"85",x"38",x"A9",x"1E",x"85", -- 0x0C20
    x"3C",x"58",x"A0",x"02",x"20",x"AB",x"AE",x"AD", -- 0x0C28
    x"A0",x"1D",x"29",x"01",x"F0",x"07",x"60",x"A0", -- 0x0C30
    x"01",x"20",x"13",x"B2",x"60",x"AD",x"A9",x"1D", -- 0x0C38
    x"C9",x"1E",x"D0",x"0C",x"A2",x"04",x"8E",x"A9", -- 0x0C40
    x"1D",x"E8",x"E8",x"8E",x"AA",x"1D",x"D0",x"15", -- 0x0C48
    x"AD",x"AA",x"1D",x"C9",x"20",x"D0",x"08",x"EE", -- 0x0C50
    x"A9",x"1D",x"EE",x"A9",x"1D",x"D0",x"06",x"EE", -- 0x0C58
    x"AA",x"1D",x"EE",x"AA",x"1D",x"AE",x"A9",x"1D", -- 0x0C60
    x"E0",x"04",x"F0",x"7E",x"CE",x"A9",x"1D",x"CE", -- 0x0C68
    x"A9",x"1D",x"AD",x"A9",x"1D",x"18",x"65",x"5E", -- 0x0C70
    x"85",x"A3",x"A5",x"5F",x"85",x"A4",x"20",x"90", -- 0x0C78
    x"B2",x"AD",x"A9",x"1D",x"0A",x"18",x"65",x"5F", -- 0x0C80
    x"85",x"A4",x"20",x"90",x"B2",x"E6",x"A4",x"20", -- 0x0C88
    x"90",x"B2",x"A5",x"5E",x"85",x"A3",x"20",x"90", -- 0x0C90
    x"B2",x"C6",x"A4",x"20",x"90",x"B2",x"A5",x"5E", -- 0x0C98
    x"38",x"ED",x"A9",x"1D",x"85",x"A3",x"20",x"90", -- 0x0CA0
    x"B2",x"E6",x"A4",x"20",x"90",x"B2",x"A5",x"5F", -- 0x0CA8
    x"85",x"A4",x"20",x"90",x"B2",x"A5",x"5F",x"38", -- 0x0CB0
    x"ED",x"A9",x"1D",x"ED",x"A9",x"1D",x"85",x"A4", -- 0x0CB8
    x"20",x"90",x"B2",x"C6",x"A4",x"20",x"90",x"B2", -- 0x0CC0
    x"A5",x"5E",x"85",x"A3",x"20",x"90",x"B2",x"E6", -- 0x0CC8
    x"A4",x"20",x"90",x"B2",x"AD",x"A9",x"1D",x"18", -- 0x0CD0
    x"65",x"5E",x"85",x"A3",x"20",x"90",x"B2",x"C6", -- 0x0CD8
    x"A4",x"20",x"90",x"B2",x"EE",x"A9",x"1D",x"EE", -- 0x0CE0
    x"A9",x"1D",x"AD",x"AA",x"1D",x"C9",x"06",x"D0", -- 0x0CE8
    x"69",x"A9",x"1E",x"18",x"65",x"5E",x"85",x"A3", -- 0x0CF0
    x"A5",x"5F",x"85",x"A4",x"20",x"90",x"B2",x"A9", -- 0x0CF8
    x"3C",x"18",x"65",x"5F",x"85",x"A4",x"20",x"90", -- 0x0D00
    x"B2",x"E6",x"A4",x"20",x"90",x"B2",x"A5",x"5E", -- 0x0D08
    x"85",x"A3",x"20",x"90",x"B2",x"C6",x"A4",x"20", -- 0x0D10
    x"90",x"B2",x"A5",x"5E",x"38",x"E9",x"1E",x"85", -- 0x0D18
    x"A3",x"20",x"90",x"B2",x"E6",x"A4",x"20",x"90", -- 0x0D20
    x"B2",x"A5",x"5F",x"85",x"A4",x"20",x"90",x"B2", -- 0x0D28
    x"A5",x"5F",x"38",x"E9",x"3C",x"85",x"A4",x"20", -- 0x0D30
    x"90",x"B2",x"C6",x"A4",x"20",x"90",x"B2",x"A5", -- 0x0D38
    x"5E",x"85",x"A3",x"20",x"90",x"B2",x"E6",x"A4", -- 0x0D40
    x"20",x"90",x"B2",x"A9",x"1E",x"18",x"65",x"5E", -- 0x0D48
    x"85",x"A3",x"20",x"90",x"B2",x"C6",x"A4",x"20", -- 0x0D50
    x"90",x"B2",x"AD",x"A9",x"1D",x"8D",x"AB",x"1D", -- 0x0D58
    x"18",x"65",x"5E",x"85",x"A3",x"A5",x"5F",x"85", -- 0x0D60
    x"A4",x"20",x"81",x"B2",x"AD",x"AB",x"1D",x"0A", -- 0x0D68
    x"18",x"65",x"5F",x"85",x"A4",x"20",x"81",x"B2", -- 0x0D70
    x"E6",x"A4",x"20",x"81",x"B2",x"A5",x"5E",x"85", -- 0x0D78
    x"A3",x"20",x"81",x"B2",x"C6",x"A4",x"20",x"81", -- 0x0D80
    x"B2",x"A5",x"5E",x"38",x"ED",x"AB",x"1D",x"85", -- 0x0D88
    x"A3",x"20",x"81",x"B2",x"E6",x"A4",x"20",x"81", -- 0x0D90
    x"B2",x"A5",x"5F",x"85",x"A4",x"20",x"81",x"B2", -- 0x0D98
    x"A5",x"5F",x"38",x"ED",x"AB",x"1D",x"ED",x"AB", -- 0x0DA0
    x"1D",x"85",x"A4",x"20",x"81",x"B2",x"C6",x"A4", -- 0x0DA8
    x"20",x"81",x"B2",x"A5",x"5E",x"85",x"A3",x"20", -- 0x0DB0
    x"81",x"B2",x"E6",x"A4",x"20",x"81",x"B2",x"AD", -- 0x0DB8
    x"AB",x"1D",x"18",x"65",x"5E",x"85",x"A3",x"20", -- 0x0DC0
    x"81",x"B2",x"C6",x"A4",x"20",x"81",x"B2",x"EE", -- 0x0DC8
    x"AB",x"1D",x"EE",x"AB",x"1D",x"AD",x"AB",x"1D", -- 0x0DD0
    x"CD",x"AA",x"1D",x"D0",x"83",x"60",x"41",x"33", -- 0x0DD8
    x"10",x"3F",x"1C",x"20",x"40",x"24",x"28",x"11", -- 0x0DE0
    x"10",x"12",x"11",x"13",x"10",x"13",x"0F",x"13", -- 0x0DE8
    x"0E",x"13",x"0D",x"12",x"0C",x"11",x"0B",x"10", -- 0x0DF0
    x"0B",x"0F",x"0C",x"0E",x"0D",x"0E",x"0E",x"0E", -- 0x0DF8
    x"0F",x"0E",x"10",x"0E",x"12",x"0E",x"14",x"0F", -- 0x0E00
    x"16",x"11",x"18",x"13",x"18",x"15",x"16",x"16", -- 0x0E08
    x"14",x"17",x"12",x"17",x"10",x"17",x"0E",x"17", -- 0x0E10
    x"0C",x"17",x"0A",x"16",x"08",x"15",x"06",x"12", -- 0x0E18
    x"04",x"0F",x"03",x"0C",x"04",x"0A",x"07",x"08", -- 0x0E20
    x"0A",x"08",x"0D",x"08",x"10",x"08",x"13",x"08", -- 0x0E28
    x"16",x"0A",x"19",x"0C",x"1C",x"0F",x"1F",x"12", -- 0x0E30
    x"20",x"15",x"20",x"00",x"03",x"06",x"FF",x"24", -- 0x0E38
    x"26",x"27",x"27",x"27",x"26",x"24",x"22",x"21", -- 0x0E40
    x"21",x"21",x"22",x"25",x"25",x"23",x"23",x"FF", -- 0x0E48
    x"51",x"53",x"55",x"58",x"5B",x"5D",x"5F",x"5D", -- 0x0E50
    x"5B",x"58",x"55",x"53",x"56",x"5A",x"5A",x"56", -- 0x0E58
    x"A9",x"00",x"8D",x"B0",x"1D",x"99",x"3C",x"03", -- 0x0E60
    x"8D",x"B1",x"1D",x"A9",x"42",x"99",x"56",x"03", -- 0x0E68
    x"AD",x"70",x"03",x"38",x"F9",x"70",x"03",x"8D", -- 0x0E70
    x"AE",x"1D",x"AD",x"8A",x"03",x"38",x"F9",x"8A", -- 0x0E78
    x"03",x"AA",x"AD",x"AE",x"1D",x"84",x"BF",x"A8", -- 0x0E80
    x"8A",x"0A",x"8A",x"6A",x"AA",x"98",x"0A",x"98", -- 0x0E88
    x"6A",x"E0",x"05",x"90",x"04",x"E0",x"FC",x"90", -- 0x0E90
    x"EE",x"C9",x"03",x"90",x"04",x"C9",x"FE",x"90", -- 0x0E98
    x"E6",x"A4",x"BF",x"8D",x"AE",x"1D",x"8A",x"8D", -- 0x0EA0
    x"AF",x"1D",x"60",x"B9",x"3C",x"03",x"30",x"2E", -- 0x0EA8
    x"B9",x"70",x"03",x"BE",x"56",x"03",x"E0",x"41", -- 0x0EB0
    x"D0",x"06",x"ED",x"AE",x"1D",x"4C",x"C7",x"AE", -- 0x0EB8
    x"E0",x"44",x"B0",x"19",x"6D",x"AE",x"1D",x"30", -- 0x0EC0
    x"15",x"C9",x"40",x"B0",x"11",x"99",x"70",x"03", -- 0x0EC8
    x"B9",x"8A",x"03",x"6D",x"AF",x"1D",x"C9",x"A0", -- 0x0ED0
    x"B0",x"04",x"99",x"8A",x"03",x"60",x"A9",x"FF", -- 0x0ED8
    x"99",x"3C",x"03",x"20",x"13",x"B2",x"60",x"20", -- 0x0EE0
    x"56",x"B0",x"A5",x"1F",x"C9",x"05",x"90",x"0F", -- 0x0EE8
    x"AD",x"14",x"91",x"CD",x"71",x"1D",x"90",x"04", -- 0x0EF0
    x"A5",x"64",x"F0",x"03",x"20",x"F5",x"A6",x"A0", -- 0x0EF8
    x"01",x"B9",x"3C",x"03",x"F0",x"22",x"A5",x"7E", -- 0x0F00
    x"18",x"69",x"10",x"99",x"70",x"03",x"A5",x"7D", -- 0x0F08
    x"18",x"69",x"16",x"99",x"8A",x"03",x"A9",x"42", -- 0x0F10
    x"99",x"56",x"03",x"20",x"60",x"AE",x"78",x"A9", -- 0x0F18
    x"51",x"85",x"36",x"A9",x"01",x"85",x"3A",x"58", -- 0x0F20
    x"A0",x"01",x"20",x"AB",x"AE",x"A0",x"02",x"20", -- 0x0F28
    x"AB",x"AE",x"AD",x"44",x"1D",x"F0",x"0D",x"A2", -- 0x0F30
    x"00",x"20",x"45",x"B7",x"A9",x"43",x"20",x"AD", -- 0x0F38
    x"B2",x"20",x"50",x"B2",x"A5",x"7E",x"C9",x"01", -- 0x0F40
    x"F0",x"16",x"C9",x"29",x"F0",x"21",x"24",x"7F", -- 0x0F48
    x"50",x"07",x"38",x"20",x"3E",x"B3",x"E6",x"7E", -- 0x0F50
    x"60",x"18",x"20",x"3E",x"B3",x"C6",x"7E",x"60", -- 0x0F58
    x"A5",x"7F",x"29",x"80",x"18",x"69",x"40",x"85", -- 0x0F60
    x"7F",x"20",x"7B",x"AF",x"4C",x"52",x"AF",x"A5", -- 0x0F68
    x"7F",x"29",x"80",x"85",x"7F",x"20",x"7B",x"AF", -- 0x0F70
    x"4C",x"59",x"AF",x"A5",x"7E",x"85",x"A3",x"C6", -- 0x0F78
    x"A3",x"A5",x"7D",x"85",x"A4",x"20",x"CD",x"AF", -- 0x0F80
    x"A5",x"7D",x"C9",x"31",x"90",x"33",x"C9",x"4F", -- 0x0F88
    x"B0",x"26",x"24",x"7F",x"10",x"11",x"A5",x"7D", -- 0x0F90
    x"85",x"A4",x"A9",x"17",x"85",x"80",x"38",x"20", -- 0x0F98
    x"E5",x"B2",x"E6",x"7D",x"E6",x"7D",x"60",x"A5", -- 0x0FA0
    x"7D",x"85",x"A4",x"A9",x"18",x"85",x"80",x"18", -- 0x0FA8
    x"20",x"E5",x"B2",x"C6",x"7D",x"C6",x"7D",x"60", -- 0x0FB0
    x"A5",x"7F",x"29",x"40",x"85",x"7F",x"4C",x"A7", -- 0x0FB8
    x"AF",x"A5",x"7F",x"29",x"40",x"18",x"69",x"80", -- 0x0FC0
    x"85",x"7F",x"4C",x"96",x"AF",x"A5",x"A3",x"85", -- 0x0FC8
    x"B3",x"A9",x"03",x"85",x"0B",x"A9",x"15",x"85", -- 0x0FD0
    x"0C",x"A5",x"B3",x"85",x"A3",x"20",x"29",x"B1", -- 0x0FD8
    x"A4",x"0B",x"A2",x"00",x"20",x"1C",x"B0",x"A5", -- 0x0FE0
    x"B3",x"18",x"69",x"10",x"85",x"A3",x"20",x"29", -- 0x0FE8
    x"B1",x"A9",x"03",x"38",x"E5",x"0B",x"A8",x"A2", -- 0x0FF0
    x"02",x"20",x"1C",x"B0",x"A4",x"0C",x"B1",x"07", -- 0x0FF8
    x"85",x"0D",x"20",x"34",x"B0",x"85",x"0E",x"B1", -- 0x1000
    x"09",x"85",x"0D",x"20",x"34",x"B0",x"91",x"07", -- 0x1008
    x"A5",x"0E",x"91",x"09",x"88",x"10",x"E7",x"C6", -- 0x1010
    x"0B",x"10",x"BA",x"60",x"B9",x"2C",x"B0",x"18", -- 0x1018
    x"65",x"A5",x"95",x"07",x"B9",x"30",x"B0",x"65", -- 0x1020
    x"A6",x"95",x"08",x"60",x"00",x"B0",x"60",x"10", -- 0x1028
    x"00",x"00",x"01",x"02",x"8D",x"73",x"03",x"A2", -- 0x1030
    x"03",x"2C",x"73",x"03",x"70",x"03",x"18",x"90", -- 0x1038
    x"01",x"38",x"66",x"0D",x"2E",x"73",x"03",x"66", -- 0x1040
    x"0D",x"2E",x"73",x"03",x"CA",x"10",x"EA",x"A5", -- 0x1048
    x"0D",x"60",x"A2",x"00",x"F0",x"02",x"A2",x"40", -- 0x1050
    x"A9",x"72",x"85",x"A4",x"86",x"72",x"A2",x"22", -- 0x1058
    x"86",x"6D",x"E8",x"E8",x"86",x"6E",x"A9",x"03", -- 0x1060
    x"85",x"6B",x"A4",x"6B",x"B9",x"D0",x"B0",x"85", -- 0x1068
    x"6F",x"85",x"70",x"B9",x"D4",x"B0",x"85",x"71", -- 0x1070
    x"A5",x"6D",x"85",x"A3",x"20",x"AC",x"B0",x"C6", -- 0x1078
    x"6D",x"C6",x"6D",x"A5",x"6E",x"85",x"A3",x"20", -- 0x1080
    x"AC",x"B0",x"E6",x"6E",x"E6",x"6E",x"C6",x"70", -- 0x1088
    x"D0",x"E6",x"24",x"72",x"70",x"04",x"E6",x"A4", -- 0x1090
    x"D0",x"02",x"C6",x"A4",x"C6",x"71",x"F0",x"07", -- 0x1098
    x"A5",x"6F",x"85",x"70",x"4C",x"78",x"B0",x"C6", -- 0x10A0
    x"6B",x"10",x"BF",x"60",x"4A",x"A8",x"29",x"07", -- 0x10A8
    x"49",x"07",x"AA",x"98",x"4A",x"4A",x"4A",x"A8", -- 0x10B0
    x"A9",x"82",x"85",x"A9",x"A9",x"BE",x"85",x"AA", -- 0x10B8
    x"BD",x"A1",x"B2",x"39",x"74",x"00",x"D0",x"04", -- 0x10C0
    x"20",x"C6",x"B1",x"60",x"20",x"0D",x"B2",x"60", -- 0x10C8
    x"01",x"02",x"03",x"02",x"04",x"03",x"02",x"01", -- 0x10D0
    x"A9",x"00",x"85",x"B1",x"85",x"B2",x"78",x"A2", -- 0x10D8
    x"7F",x"8E",x"22",x"91",x"AD",x"20",x"91",x"29", -- 0x10E0
    x"80",x"D0",x"02",x"E6",x"B1",x"A2",x"FF",x"8E", -- 0x10E8
    x"22",x"91",x"A2",x"F7",x"8E",x"20",x"91",x"58", -- 0x10F0
    x"AD",x"11",x"91",x"CD",x"11",x"91",x"D0",x"F8", -- 0x10F8
    x"A2",x"00",x"29",x"3E",x"C9",x"1F",x"B0",x"06", -- 0x1100
    x"A6",x"B0",x"D0",x"02",x"A2",x"80",x"86",x"B0", -- 0x1108
    x"29",x"1F",x"C9",x"0F",x"B0",x"02",x"C6",x"B1", -- 0x1110
    x"A2",x"02",x"29",x"0F",x"C9",x"08",x"90",x"06", -- 0x1118
    x"A2",x"FE",x"29",x"04",x"D0",x"02",x"86",x"B2", -- 0x1120
    x"60",x"A5",x"A4",x"C9",x"B0",x"B0",x"2D",x"A5", -- 0x1128
    x"A3",x"C9",x"48",x"B0",x"27",x"29",x"03",x"85", -- 0x1130
    x"AD",x"A5",x"A3",x"4A",x"29",x"FE",x"AA",x"18", -- 0x1138
    x"BD",x"5F",x"B1",x"65",x"A4",x"85",x"A5",x"BD", -- 0x1140
    x"60",x"B1",x"69",x"00",x"85",x"A6",x"18",x"A5", -- 0x1148
    x"A5",x"69",x"B0",x"85",x"A7",x"A5",x"A6",x"69", -- 0x1150
    x"00",x"85",x"A8",x"60",x"68",x"68",x"60",x"00", -- 0x1158
    x"10",x"B0",x"10",x"60",x"11",x"10",x"12",x"C0", -- 0x1160
    x"12",x"70",x"13",x"20",x"14",x"D0",x"14",x"80", -- 0x1168
    x"15",x"30",x"16",x"E0",x"16",x"90",x"17",x"40", -- 0x1170
    x"18",x"F0",x"18",x"A0",x"19",x"50",x"1A",x"00", -- 0x1178
    x"1B",x"B0",x"1B",x"20",x"29",x"B1",x"4C",x"CD", -- 0x1180
    x"B1",x"B9",x"56",x"03",x"AA",x"20",x"AD",x"B2", -- 0x1188
    x"B9",x"70",x"03",x"85",x"A3",x"B9",x"8A",x"03", -- 0x1190
    x"85",x"A4",x"8A",x"C9",x"38",x"90",x"04",x"C9", -- 0x1198
    x"46",x"90",x"23",x"20",x"BB",x"B1",x"A5",x"A3", -- 0x11A0
    x"18",x"69",x"04",x"85",x"A3",x"18",x"A9",x"10", -- 0x11A8
    x"65",x"A9",x"85",x"A9",x"90",x"02",x"E6",x"AA", -- 0x11B0
    x"4C",x"BF",x"B1",x"A9",x"00",x"85",x"1A",x"20", -- 0x11B8
    x"29",x"B1",x"A0",x"0F",x"D0",x"09",x"A9",x"00", -- 0x11C0
    x"85",x"1A",x"20",x"29",x"B1",x"A0",x"07",x"B1", -- 0x11C8
    x"A9",x"A2",x"00",x"86",x"AC",x"A6",x"AD",x"F0", -- 0x11D0
    x"0A",x"18",x"4A",x"66",x"AC",x"4A",x"66",x"AC", -- 0x11D8
    x"CA",x"D0",x"F7",x"85",x"AB",x"B1",x"A5",x"F0", -- 0x11E0
    x"08",x"AA",x"25",x"AB",x"05",x"1A",x"85",x"1A", -- 0x11E8
    x"8A",x"05",x"AB",x"91",x"A5",x"A5",x"AD",x"F0", -- 0x11F0
    x"10",x"B1",x"A7",x"F0",x"08",x"AA",x"25",x"AC", -- 0x11F8
    x"05",x"1A",x"85",x"1A",x"8A",x"05",x"AC",x"91", -- 0x1200
    x"A7",x"88",x"10",x"C3",x"60",x"20",x"29",x"B1", -- 0x1208
    x"4C",x"57",x"B2",x"B9",x"56",x"03",x"AA",x"20", -- 0x1210
    x"AD",x"B2",x"B9",x"A4",x"03",x"85",x"A3",x"B9", -- 0x1218
    x"BE",x"03",x"85",x"A4",x"8A",x"C9",x"38",x"90", -- 0x1220
    x"04",x"C9",x"46",x"90",x"23",x"20",x"45",x"B2", -- 0x1228
    x"A5",x"A3",x"18",x"69",x"04",x"85",x"A3",x"18", -- 0x1230
    x"A9",x"10",x"65",x"A9",x"85",x"A9",x"90",x"02", -- 0x1238
    x"E6",x"AA",x"4C",x"49",x"B2",x"A9",x"00",x"85", -- 0x1240
    x"1A",x"20",x"29",x"B1",x"A0",x"0F",x"D0",x"09", -- 0x1248
    x"A9",x"00",x"85",x"1A",x"20",x"29",x"B1",x"A0", -- 0x1250
    x"07",x"B1",x"A9",x"49",x"FF",x"A2",x"FF",x"86", -- 0x1258
    x"AC",x"A6",x"AD",x"F0",x"0A",x"38",x"6A",x"66", -- 0x1260
    x"AC",x"6A",x"66",x"AC",x"CA",x"D0",x"F7",x"31", -- 0x1268
    x"A5",x"91",x"A5",x"A5",x"AD",x"F0",x"06",x"A5", -- 0x1270
    x"AC",x"31",x"A7",x"91",x"A7",x"88",x"10",x"D9", -- 0x1278
    x"60",x"20",x"29",x"B1",x"A6",x"AD",x"BD",x"A9", -- 0x1280
    x"B2",x"A2",x"00",x"01",x"A5",x"81",x"A5",x"60", -- 0x1288
    x"20",x"29",x"B1",x"A6",x"AD",x"BD",x"A9",x"B2", -- 0x1290
    x"A2",x"00",x"49",x"FF",x"21",x"A5",x"81",x"A5", -- 0x1298
    x"60",x"80",x"40",x"20",x"10",x"08",x"04",x"02", -- 0x12A0
    x"01",x"C0",x"30",x"0C",x"03",x"85",x"29",x"A9", -- 0x12A8
    x"00",x"85",x"AA",x"A5",x"29",x"0A",x"26",x"AA", -- 0x12B0
    x"0A",x"26",x"AA",x"0A",x"26",x"AA",x"18",x"69", -- 0x12B8
    x"02",x"85",x"A9",x"A5",x"AA",x"69",x"BB",x"85", -- 0x12C0
    x"AA",x"60",x"85",x"29",x"A9",x"00",x"85",x"AA", -- 0x12C8
    x"A5",x"29",x"0A",x"26",x"AA",x"0A",x"26",x"AA", -- 0x12D0
    x"0A",x"26",x"AA",x"85",x"A9",x"A5",x"AA",x"18", -- 0x12D8
    x"69",x"80",x"85",x"AA",x"60",x"C6",x"A4",x"C6", -- 0x12E0
    x"A4",x"A9",x"11",x"85",x"58",x"B0",x"13",x"20", -- 0x12E8
    x"13",x"B3",x"A0",x"00",x"B1",x"A7",x"91",x"A5", -- 0x12F0
    x"C8",x"C4",x"80",x"D0",x"F7",x"C6",x"58",x"10", -- 0x12F8
    x"EE",x"60",x"20",x"13",x"B3",x"A4",x"80",x"B1", -- 0x1300
    x"A5",x"91",x"A7",x"88",x"10",x"F9",x"C6",x"58", -- 0x1308
    x"10",x"F0",x"60",x"A6",x"58",x"BD",x"2B",x"B3", -- 0x1310
    x"85",x"A3",x"20",x"29",x"B1",x"18",x"A5",x"A5", -- 0x1318
    x"69",x"02",x"85",x"A7",x"A5",x"A6",x"69",x"00", -- 0x1320
    x"85",x"A8",x"60",x"00",x"04",x"08",x"0C",x"10", -- 0x1328
    x"14",x"18",x"1C",x"20",x"24",x"28",x"2C",x"30", -- 0x1330
    x"34",x"38",x"3C",x"40",x"44",x"48",x"A0",x"15", -- 0x1338
    x"B0",x"3E",x"84",x"80",x"A5",x"7E",x"18",x"69", -- 0x1340
    x"1E",x"85",x"A3",x"A5",x"7D",x"85",x"A4",x"20", -- 0x1348
    x"29",x"B1",x"A4",x"80",x"A9",x"00",x"85",x"0E", -- 0x1350
    x"A9",x"09",x"85",x"0F",x"18",x"66",x"0E",x"66", -- 0x1358
    x"0E",x"B1",x"A5",x"2A",x"26",x"0E",x"2A",x"91", -- 0x1360
    x"A5",x"26",x"0E",x"A5",x"A5",x"38",x"E9",x"B0", -- 0x1368
    x"85",x"A5",x"A5",x"A6",x"E9",x"00",x"85",x"A6", -- 0x1370
    x"C6",x"0F",x"D0",x"E0",x"88",x"10",x"C3",x"60", -- 0x1378
    x"84",x"80",x"A5",x"7E",x"85",x"A3",x"A5",x"7D", -- 0x1380
    x"85",x"A4",x"20",x"29",x"B1",x"A4",x"80",x"A9", -- 0x1388
    x"00",x"85",x"0E",x"A9",x"09",x"85",x"0F",x"18", -- 0x1390
    x"26",x"0E",x"26",x"0E",x"B1",x"A5",x"6A",x"66", -- 0x1398
    x"0E",x"6A",x"91",x"A5",x"66",x"0E",x"A5",x"A5", -- 0x13A0
    x"18",x"69",x"B0",x"85",x"A5",x"A5",x"A6",x"69", -- 0x13A8
    x"00",x"85",x"A6",x"C6",x"0F",x"D0",x"E0",x"88", -- 0x13B0
    x"10",x"C6",x"60",x"20",x"DF",x"A3",x"A9",x"FF", -- 0x13B8
    x"A2",x"18",x"9D",x"3C",x"03",x"CA",x"10",x"FA", -- 0x13C0
    x"E8",x"86",x"64",x"8E",x"6F",x"03",x"AD",x"0E", -- 0x13C8
    x"90",x"29",x"0F",x"09",x"10",x"8D",x"0E",x"90", -- 0x13D0
    x"A9",x"6A",x"8D",x"0F",x"90",x"A9",x"01",x"A2", -- 0x13D8
    x"90",x"9D",x"35",x"96",x"CA",x"D0",x"FA",x"78", -- 0x13E0
    x"F8",x"A5",x"81",x"18",x"69",x"01",x"85",x"81", -- 0x13E8
    x"D8",x"58",x"20",x"08",x"B4",x"A9",x"48",x"85", -- 0x13F0
    x"BE",x"20",x"F5",x"A6",x"20",x"A6",x"A4",x"A9", -- 0x13F8
    x"15",x"20",x"96",x"B9",x"C6",x"BE",x"D0",x"F1", -- 0x1400
    x"A9",x"0A",x"85",x"A3",x"A9",x"30",x"85",x"A4", -- 0x1408
    x"A0",x"00",x"B9",x"32",x"B6",x"20",x"81",x"B5", -- 0x1410
    x"C0",x"05",x"D0",x"F6",x"A5",x"1F",x"C9",x"14", -- 0x1418
    x"90",x"04",x"A0",x"05",x"B0",x"05",x"4A",x"4A", -- 0x1420
    x"29",x"07",x"A8",x"A9",x"22",x"85",x"A3",x"B9", -- 0x1428
    x"D7",x"B5",x"A8",x"18",x"69",x"07",x"85",x"80", -- 0x1430
    x"B9",x"DD",x"B5",x"20",x"81",x"B5",x"C4",x"80", -- 0x1438
    x"D0",x"F6",x"A9",x"0E",x"85",x"A3",x"A9",x"58", -- 0x1440
    x"85",x"A4",x"A0",x"00",x"84",x"B3",x"B9",x"07", -- 0x1448
    x"B6",x"20",x"81",x"B5",x"C0",x"08",x"D0",x"F6", -- 0x1450
    x"A9",x"32",x"85",x"A3",x"A5",x"81",x"29",x"F0", -- 0x1458
    x"4A",x"4A",x"4A",x"4A",x"20",x"51",x"B5",x"A9", -- 0x1460
    x"36",x"85",x"A3",x"A9",x"FF",x"85",x"72",x"A5", -- 0x1468
    x"81",x"29",x"0F",x"20",x"51",x"B5",x"A5",x"1F", -- 0x1470
    x"29",x"03",x"A8",x"B9",x"0F",x"B6",x"A8",x"B9", -- 0x1478
    x"13",x"B6",x"85",x"A3",x"A9",x"78",x"85",x"A4", -- 0x1480
    x"C8",x"84",x"80",x"B9",x"13",x"B6",x"18",x"65", -- 0x1488
    x"80",x"85",x"80",x"C8",x"B9",x"13",x"B6",x"20", -- 0x1490
    x"81",x"B5",x"C4",x"80",x"D0",x"F6",x"A9",x"00", -- 0x1498
    x"85",x"A3",x"A8",x"A9",x"A0",x"85",x"A4",x"B9", -- 0x14A0
    x"47",x"B6",x"20",x"81",x"B5",x"C0",x"0B",x"D0", -- 0x14A8
    x"F6",x"A9",x"30",x"85",x"A3",x"A2",x"02",x"B5", -- 0x14B0
    x"22",x"95",x"1B",x"CA",x"10",x"F9",x"20",x"2E", -- 0x14B8
    x"B5",x"20",x"F2",x"B4",x"A9",x"00",x"85",x"A3", -- 0x14C0
    x"85",x"A4",x"A0",x"60",x"84",x"B3",x"98",x"20", -- 0x14C8
    x"AD",x"B2",x"20",x"86",x"B5",x"C0",x"65",x"D0", -- 0x14D0
    x"F3",x"F0",x"06",x"A9",x"00",x"85",x"72",x"85", -- 0x14D8
    x"A4",x"A9",x"14",x"85",x"A3",x"A2",x"02",x"B5", -- 0x14E0
    x"F7",x"95",x"1B",x"CA",x"10",x"F9",x"20",x"2E", -- 0x14E8
    x"B5",x"60",x"A9",x"30",x"85",x"A3",x"A2",x"00", -- 0x14F0
    x"86",x"A4",x"86",x"80",x"A9",x"A0",x"20",x"CA", -- 0x14F8
    x"B2",x"20",x"0D",x"B2",x"20",x"77",x"B5",x"E8", -- 0x1500
    x"E0",x"06",x"D0",x"EE",x"A5",x"1E",x"F0",x"1D", -- 0x1508
    x"85",x"80",x"C6",x"80",x"F0",x"17",x"A9",x"44", -- 0x1510
    x"85",x"A3",x"A9",x"6F",x"20",x"AD",x"B2",x"20", -- 0x1518
    x"C6",x"B1",x"A5",x"A3",x"38",x"E9",x"04",x"85", -- 0x1520
    x"A3",x"C6",x"80",x"D0",x"ED",x"60",x"A2",x"02", -- 0x1528
    x"A9",x"00",x"85",x"72",x"F0",x"0B",x"B5",x"1B", -- 0x1530
    x"29",x"F0",x"4A",x"4A",x"4A",x"4A",x"20",x"51", -- 0x1538
    x"B5",x"B5",x"1B",x"29",x"0F",x"20",x"51",x"B5", -- 0x1540
    x"CA",x"10",x"EB",x"A9",x"00",x"20",x"51",x"B5", -- 0x1548
    x"60",x"85",x"0E",x"86",x"80",x"A9",x"A0",x"20", -- 0x1550
    x"CA",x"B2",x"20",x"0D",x"B2",x"A5",x"0E",x"F0", -- 0x1558
    x"07",x"A9",x"FF",x"85",x"72",x"4C",x"6C",x"B5", -- 0x1560
    x"24",x"72",x"10",x"0B",x"A5",x"0E",x"18",x"69", -- 0x1568
    x"65",x"20",x"AD",x"B2",x"20",x"C6",x"B1",x"A5", -- 0x1570
    x"A3",x"18",x"69",x"04",x"85",x"A3",x"A6",x"80", -- 0x1578
    x"60",x"84",x"B3",x"20",x"CA",x"B2",x"20",x"C6", -- 0x1580
    x"B1",x"A5",x"A3",x"18",x"69",x"04",x"85",x"A3", -- 0x1588
    x"A4",x"B3",x"C8",x"60",x"20",x"BB",x"B3",x"A9", -- 0x1590
    x"0A",x"85",x"A3",x"A9",x"78",x"85",x"A4",x"A9", -- 0x1598
    x"A0",x"20",x"CA",x"B2",x"A0",x"0E",x"84",x"B3", -- 0x15A0
    x"20",x"0D",x"B2",x"A5",x"A3",x"18",x"69",x"04", -- 0x15A8
    x"85",x"A3",x"C6",x"B3",x"D0",x"F2",x"A9",x"0A", -- 0x15B0
    x"85",x"A3",x"A0",x"00",x"B9",x"CA",x"B5",x"20", -- 0x15B8
    x"81",x"B5",x"C0",x"0D",x"D0",x"F6",x"20",x"8E", -- 0x15C0
    x"B9",x"60",x"02",x"09",x"14",x"05",x"20",x"14", -- 0x15C8
    x"08",x"05",x"20",x"04",x"15",x"13",x"14",x"00", -- 0x15D0
    x"07",x"0E",x"15",x"1C",x"23",x"20",x"03",x"01", -- 0x15D8
    x"04",x"05",x"14",x"20",x"03",x"01",x"10",x"14", -- 0x15E0
    x"01",x"09",x"0E",x"03",x"0F",x"0C",x"0F",x"0E", -- 0x15E8
    x"05",x"0C",x"07",x"05",x"0E",x"05",x"12",x"01", -- 0x15F0
    x"0C",x"17",x"01",x"12",x"12",x"09",x"0F",x"12", -- 0x15F8
    x"01",x"16",x"05",x"0E",x"07",x"05",x"12",x"0D", -- 0x1600
    x"09",x"13",x"13",x"09",x"0F",x"0E",x"3A",x"00", -- 0x1608
    x"0F",x"1D",x"29",x"0A",x"0E",x"01",x"13",x"14", -- 0x1610
    x"12",x"0F",x"20",x"02",x"01",x"14",x"14",x"0C", -- 0x1618
    x"05",x"13",x"0C",x"0D",x"0C",x"01",x"13",x"05", -- 0x1620
    x"12",x"20",x"01",x"14",x"14",x"01",x"03",x"0B", -- 0x1628
    x"10",x"0B",x"13",x"10",x"01",x"03",x"05",x"20", -- 0x1630
    x"17",x"01",x"12",x"10",x"12",x"0A",x"06",x"0C", -- 0x1638
    x"01",x"07",x"20",x"13",x"08",x"09",x"10",x"08", -- 0x1640
    x"09",x"07",x"08",x"20",x"13",x"03",x"0F",x"12", -- 0x1648
    x"05",x"3A",x"A2",x"00",x"86",x"AE",x"20",x"45", -- 0x1650
    x"B7",x"A9",x"43",x"20",x"AD",x"B2",x"20",x"50", -- 0x1658
    x"B2",x"78",x"A9",x"07",x"85",x"37",x"85",x"38", -- 0x1660
    x"A9",x"01",x"85",x"3B",x"85",x"3C",x"58",x"85", -- 0x1668
    x"B0",x"AD",x"70",x"03",x"18",x"69",x"03",x"8D", -- 0x1670
    x"4A",x"1D",x"A9",x"F9",x"8D",x"3E",x"1D",x"AD", -- 0x1678
    x"8A",x"03",x"18",x"69",x"FE",x"8D",x"50",x"1D", -- 0x1680
    x"A9",x"96",x"8D",x"44",x"1D",x"A9",x"00",x"8D", -- 0x1688
    x"56",x"1D",x"60",x"A9",x"00",x"85",x"1A",x"85", -- 0x1690
    x"25",x"85",x"AE",x"A9",x"05",x"85",x"B4",x"A6", -- 0x1698
    x"B4",x"BD",x"44",x"1D",x"F0",x"5B",x"20",x"45", -- 0x16A0
    x"B7",x"A9",x"43",x"20",x"AD",x"B2",x"20",x"50", -- 0x16A8
    x"B2",x"A6",x"B4",x"DE",x"44",x"1D",x"F0",x"74", -- 0x16B0
    x"BD",x"4A",x"1D",x"85",x"A3",x"A5",x"20",x"C9", -- 0x16B8
    x"03",x"D0",x"23",x"A5",x"7D",x"CD",x"50",x"1D", -- 0x16C0
    x"B0",x"1C",x"69",x"16",x"CD",x"50",x"1D",x"90", -- 0x16C8
    x"15",x"A5",x"7E",x"CD",x"4A",x"1D",x"F0",x"09", -- 0x16D0
    x"B0",x"0C",x"69",x"20",x"CD",x"4A",x"1D",x"90", -- 0x16D8
    x"05",x"18",x"A9",x"FE",x"D0",x"04",x"18",x"BD", -- 0x16E0
    x"3E",x"1D",x"85",x"AF",x"7D",x"50",x"1D",x"C9", -- 0x16E8
    x"09",x"90",x"2C",x"C9",x"A8",x"B0",x"28",x"85", -- 0x16F0
    x"A4",x"9D",x"50",x"1D",x"20",x"C6",x"B1",x"A5", -- 0x16F8
    x"1A",x"F0",x"3A",x"A5",x"20",x"F0",x"0F",x"C9", -- 0x1700
    x"03",x"D0",x"32",x"A6",x"B4",x"D0",x"2E",x"20", -- 0x1708
    x"81",x"B7",x"F0",x"0B",x"D0",x"2E",x"A6",x"B4", -- 0x1710
    x"F0",x"2A",x"20",x"81",x"B7",x"D0",x"1E",x"A6", -- 0x1718
    x"B4",x"20",x"45",x"B7",x"A9",x"43",x"20",x"AD", -- 0x1720
    x"B2",x"20",x"50",x"B2",x"A6",x"B4",x"A9",x"00", -- 0x1728
    x"9D",x"44",x"1D",x"85",x"1A",x"A9",x"FF",x"9D", -- 0x1730
    x"4A",x"1D",x"9D",x"50",x"1D",x"C6",x"B4",x"30", -- 0x1738
    x"03",x"4C",x"9F",x"B6",x"60",x"BD",x"4A",x"1D", -- 0x1740
    x"85",x"A3",x"BD",x"50",x"1D",x"85",x"A4",x"BD", -- 0x1748
    x"3E",x"1D",x"85",x"AF",x"60",x"A0",x"05",x"A6", -- 0x1750
    x"2F",x"B9",x"44",x"1D",x"D0",x"1F",x"BD",x"70", -- 0x1758
    x"03",x"69",x"02",x"99",x"4A",x"1D",x"A9",x"05", -- 0x1760
    x"99",x"3E",x"1D",x"18",x"7D",x"8A",x"03",x"99", -- 0x1768
    x"50",x"1D",x"A9",x"23",x"99",x"44",x"1D",x"A9", -- 0x1770
    x"01",x"99",x"56",x"1D",x"60",x"88",x"D0",x"D9", -- 0x1778
    x"60",x"A4",x"A4",x"C9",x"00",x"F0",x"0A",x"C0", -- 0x1780
    x"67",x"90",x"2E",x"C0",x"73",x"90",x"0D",x"B0", -- 0x1788
    x"08",x"C0",x"6E",x"90",x"04",x"C0",x"7E",x"90", -- 0x1790
    x"03",x"A0",x"FF",x"60",x"A5",x"A3",x"4A",x"A8", -- 0x1798
    x"29",x"07",x"49",x"07",x"AA",x"98",x"4A",x"4A", -- 0x17A0
    x"4A",x"A8",x"BD",x"A1",x"B2",x"19",x"74",x"00", -- 0x17A8
    x"99",x"74",x"00",x"A9",x"00",x"60",x"A0",x"FF", -- 0x17B0
    x"60",x"AD",x"50",x"1D",x"C5",x"7D",x"90",x"F6", -- 0x17B8
    x"A5",x"7E",x"CD",x"4A",x"1D",x"F0",x"09",x"B0", -- 0x17C0
    x"ED",x"69",x"20",x"CD",x"4A",x"1D",x"90",x"E6", -- 0x17C8
    x"A5",x"7D",x"18",x"69",x"06",x"C5",x"A4",x"B0", -- 0x17D0
    x"7E",x"69",x"04",x"C5",x"A4",x"90",x"78",x"A5", -- 0x17D8
    x"7E",x"69",x"0A",x"C5",x"A3",x"B0",x"70",x"69", -- 0x17E0
    x"04",x"C5",x"A3",x"90",x"6A",x"78",x"A9",x"68", -- 0x17E8
    x"85",x"36",x"A9",x"02",x"85",x"3A",x"A9",x"82", -- 0x17F0
    x"85",x"38",x"A9",x"0A",x"85",x"3C",x"A9",x"04", -- 0x17F8
    x"85",x"35",x"A9",x"0A",x"85",x"39",x"F8",x"A9", -- 0x1800
    x"01",x"18",x"20",x"60",x"B9",x"A9",x"04",x"8D", -- 0x1808
    x"A9",x"1D",x"A9",x"20",x"8D",x"AA",x"1D",x"A9", -- 0x1810
    x"0C",x"85",x"B4",x"A5",x"7E",x"18",x"69",x"0E", -- 0x1818
    x"85",x"5E",x"A5",x"7D",x"18",x"69",x"0A",x"85", -- 0x1820
    x"5F",x"AD",x"0F",x"90",x"85",x"B3",x"20",x"3D", -- 0x1828
    x"AC",x"A5",x"B4",x"0A",x"0A",x"0A",x"0A",x"05", -- 0x1830
    x"B4",x"8D",x"0F",x"90",x"20",x"94",x"B9",x"C6", -- 0x1838
    x"B4",x"D0",x"EB",x"A5",x"B3",x"8D",x"0F",x"90", -- 0x1840
    x"A9",x"00",x"85",x"31",x"A5",x"1F",x"C9",x"04", -- 0x1848
    x"D0",x"4E",x"E6",x"1E",x"4C",x"A0",x"B8",x"A5", -- 0x1850
    x"7D",x"18",x"69",x"18",x"C5",x"A4",x"90",x"40", -- 0x1858
    x"A5",x"A4",x"69",x"07",x"C5",x"7D",x"90",x"38", -- 0x1860
    x"78",x"A9",x"20",x"85",x"37",x"A9",x"01",x"85", -- 0x1868
    x"3B",x"58",x"A9",x"05",x"20",x"55",x"B9",x"AD", -- 0x1870
    x"58",x"03",x"C9",x"44",x"D0",x"07",x"C9",x"45", -- 0x1878
    x"D0",x"03",x"A9",x"00",x"60",x"AD",x"4A",x"1D", -- 0x1880
    x"8D",x"72",x"03",x"A5",x"7D",x"18",x"69",x"18", -- 0x1888
    x"8D",x"8C",x"03",x"A9",x"41",x"8D",x"58",x"03", -- 0x1890
    x"A9",x"00",x"8D",x"3E",x"03",x"8D",x"28",x"1D", -- 0x1898
    x"60",x"84",x"BF",x"20",x"13",x"B2",x"A4",x"BF", -- 0x18A0
    x"B9",x"56",x"03",x"C9",x"38",x"90",x"44",x"C9", -- 0x18A8
    x"46",x"B0",x"4B",x"E9",x"37",x"AA",x"BD",x"72", -- 0x18B0
    x"B9",x"20",x"44",x"B9",x"A4",x"BF",x"B9",x"24", -- 0x18B8
    x"1D",x"D0",x"22",x"78",x"A9",x"30",x"85",x"37", -- 0x18C0
    x"A9",x"01",x"85",x"3B",x"A9",x"02",x"85",x"38", -- 0x18C8
    x"A9",x"01",x"85",x"3C",x"58",x"B9",x"A4",x"03", -- 0x18D0
    x"99",x"70",x"03",x"B9",x"BE",x"03",x"99",x"8A", -- 0x18D8
    x"03",x"A9",x"45",x"D0",x"56",x"C9",x"08",x"D0", -- 0x18E0
    x"04",x"A9",x"44",x"D0",x"4E",x"C9",x"10",x"D0", -- 0x18E8
    x"4D",x"F0",x"3E",x"4A",x"4A",x"AA",x"BD",x"80", -- 0x18F0
    x"B9",x"20",x"44",x"B9",x"A4",x"BF",x"B9",x"24", -- 0x18F8
    x"1D",x"D0",x"22",x"78",x"A9",x"04",x"85",x"35", -- 0x1900
    x"A9",x"01",x"85",x"39",x"A9",x"82",x"85",x"38", -- 0x1908
    x"A9",x"01",x"85",x"3C",x"58",x"B9",x"A4",x"03", -- 0x1910
    x"99",x"70",x"03",x"B9",x"BE",x"03",x"99",x"8A", -- 0x1918
    x"03",x"A9",x"4A",x"D0",x"16",x"C9",x"08",x"D0", -- 0x1920
    x"04",x"A9",x"46",x"D0",x"0E",x"C9",x"10",x"D0", -- 0x1928
    x"0D",x"A9",x"FF",x"99",x"3C",x"03",x"99",x"24", -- 0x1930
    x"1D",x"A9",x"35",x"99",x"56",x"03",x"A6",x"BF", -- 0x1938
    x"FE",x"24",x"1D",x"60",x"30",x"02",x"C6",x"31", -- 0x1940
    x"C9",x"FF",x"D0",x"07",x"C6",x"1E",x"85",x"3E", -- 0x1948
    x"4C",x"6C",x"B9",x"29",x"7F",x"78",x"F8",x"18", -- 0x1950
    x"65",x"F7",x"85",x"F7",x"90",x"0E",x"A9",x"00", -- 0x1958
    x"65",x"F8",x"85",x"F8",x"90",x"06",x"A9",x"00", -- 0x1960
    x"65",x"F9",x"85",x"F9",x"D8",x"58",x"20",x"DB", -- 0x1968
    x"B4",x"60",x"80",x"10",x"08",x"06",x"06",x"08", -- 0x1970
    x"10",x"10",x"10",x"10",x"80",x"80",x"80",x"80", -- 0x1978
    x"FF",x"A5",x"30",x"10",x"10",x"80",x"80",x"90", -- 0x1980
    x"90",x"90",x"90",x"A0",x"90",x"90",x"A9",x"FF", -- 0x1988
    x"85",x"19",x"D0",x"04",x"A9",x"40",x"85",x"19", -- 0x1990
    x"A9",x"FF",x"85",x"30",x"C6",x"30",x"D0",x"FC", -- 0x1998
    x"C6",x"19",x"D0",x"F4",x"60",x"A9",x"0E",x"8D", -- 0x19A0
    x"0F",x"90",x"20",x"DF",x"A3",x"A9",x"02",x"A2", -- 0x19A8
    x"C6",x"9D",x"FF",x"95",x"CA",x"D0",x"FA",x"A9", -- 0x19B0
    x"2E",x"85",x"A4",x"A2",x"09",x"A5",x"A4",x"18", -- 0x19B8
    x"69",x"08",x"85",x"A4",x"A9",x"07",x"85",x"A3", -- 0x19C0
    x"86",x"5E",x"A6",x"5E",x"BD",x"1C",x"BA",x"85", -- 0x19C8
    x"5F",x"A0",x"00",x"A5",x"5F",x"0A",x"85",x"5F", -- 0x19D0
    x"A9",x"20",x"90",x"02",x"A9",x"A0",x"20",x"81", -- 0x19D8
    x"B5",x"C0",x"08",x"D0",x"EE",x"A6",x"5E",x"CA", -- 0x19E0
    x"30",x"06",x"8A",x"4A",x"90",x"DA",x"B0",x"CD", -- 0x19E8
    x"A9",x"78",x"85",x"A4",x"A0",x"00",x"84",x"A3", -- 0x19F0
    x"B9",x"26",x"BA",x"F0",x"08",x"30",x"14",x"20", -- 0x19F8
    x"81",x"B5",x"4C",x"F8",x"B9",x"A5",x"A4",x"18", -- 0x1A00
    x"69",x"0E",x"85",x"A4",x"C8",x"A9",x"00",x"85", -- 0x1A08
    x"A3",x"F0",x"E5",x"A2",x"02",x"20",x"8E",x"B9", -- 0x1A10
    x"CA",x"10",x"FA",x"60",x"A8",x"EE",x"A8",x"AA", -- 0x1A18
    x"CC",x"8A",x"A8",x"8A",x"EE",x"EE",x"28",x"03", -- 0x1A20
    x"29",x"20",x"31",x"39",x"38",x"32",x"00",x"20", -- 0x1A28
    x"20",x"20",x"03",x"0F",x"0D",x"0D",x"0F",x"04", -- 0x1A30
    x"0F",x"12",x"05",x"20",x"0C",x"14",x"04",x"2E", -- 0x1A38
    x"00",x"28",x"03",x"29",x"20",x"31",x"39",x"38", -- 0x1A40
    x"31",x"00",x"20",x"20",x"20",x"02",x"01",x"0C", -- 0x1A48
    x"0C",x"19",x"20",x"0D",x"09",x"04",x"17",x"01", -- 0x1A50
    x"19",x"FF",x"20",x"A5",x"B9",x"AD",x"08",x"90", -- 0x1A58
    x"C9",x"02",x"B0",x"0A",x"AD",x"09",x"90",x"C9", -- 0x1A60
    x"08",x"B0",x"03",x"20",x"BB",x"BA",x"20",x"D8", -- 0x1A68
    x"B0",x"A5",x"B1",x"F0",x"0D",x"30",x"0B",x"AD", -- 0x1A70
    x"00",x"90",x"18",x"69",x"01",x"29",x"8F",x"8D", -- 0x1A78
    x"00",x"90",x"A5",x"B2",x"F0",x"0F",x"30",x"0D", -- 0x1A80
    x"AD",x"01",x"90",x"18",x"69",x"01",x"29",x"1F", -- 0x1A88
    x"8D",x"01",x"90",x"90",x"0A",x"F0",x"08",x"AD", -- 0x1A90
    x"00",x"90",x"49",x"80",x"8D",x"00",x"90",x"A5", -- 0x1A98
    x"B0",x"F0",x"12",x"A9",x"06",x"85",x"1E",x"A2", -- 0x1AA0
    x"00",x"86",x"1F",x"E8",x"86",x"42",x"86",x"81", -- 0x1AA8
    x"68",x"68",x"4C",x"2F",x"A0",x"A9",x"05",x"20", -- 0x1AB0
    x"96",x"B9",x"60",x"20",x"DF",x"A3",x"A9",x"03", -- 0x1AB8
    x"A2",x"C6",x"9D",x"FF",x"95",x"CA",x"D0",x"FA", -- 0x1AC0
    x"A9",x"0A",x"85",x"A3",x"A9",x"28",x"85",x"A4", -- 0x1AC8
    x"A0",x"00",x"B9",x"B0",x"BF",x"F0",x"08",x"30", -- 0x1AD0
    x"14",x"20",x"81",x"B5",x"4C",x"D2",x"BA",x"C8", -- 0x1AD8
    x"A5",x"A4",x"18",x"69",x"0E",x"85",x"A4",x"A9", -- 0x1AE0
    x"0A",x"85",x"A3",x"D0",x"E5",x"A9",x"0A",x"85", -- 0x1AE8
    x"BE",x"20",x"8E",x"B9",x"C6",x"BE",x"D0",x"F9", -- 0x1AF0
    x"60",x"2C",x"11",x"91",x"68",x"A8",x"68",x"AA", -- 0x1AF8
    x"68",x"40",x"01",x"05",x"05",x"01",x"81",x"85", -- 0x1B00
    x"46",x"65",x"66",x"45",x"46",x"45",x"41",x"40", -- 0x1B08
    x"C0",x"00",x"00",x"40",x"40",x"00",x"08",x"48", -- 0x1B10
    x"44",x"64",x"64",x"44",x"44",x"44",x"04",x"04", -- 0x1B18
    x"0C",x"00",x"81",x"25",x"05",x"15",x"15",x"19", -- 0x1B20
    x"19",x"15",x"15",x"1A",x"1A",x"15",x"05",x"08", -- 0x1B28
    x"08",x"28",x"08",x"60",x"40",x"50",x"50",x"90", -- 0x1B30
    x"90",x"50",x"50",x"90",x"90",x"50",x"40",x"80", -- 0x1B38
    x"80",x"A0",x"00",x"F0",x"30",x"30",x"31",x"35", -- 0x1B40
    x"35",x"35",x"05",x"05",x"02",x"02",x"02",x"02", -- 0x1B48
    x"00",x"00",x"00",x"3C",x"30",x"30",x"30",x"70", -- 0x1B50
    x"70",x"70",x"40",x"40",x"00",x"00",x"00",x"00", -- 0x1B58
    x"00",x"00",x"00",x"00",x"00",x"00",x"A0",x"20", -- 0x1B60
    x"28",x"05",x"05",x"03",x"03",x"00",x"00",x"00", -- 0x1B68
    x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"20", -- 0x1B70
    x"A0",x"40",x"40",x"00",x"00",x"00",x"00",x"00", -- 0x1B78
    x"00",x"00",x"83",x"2F",x"0F",x"3F",x"3B",x"3B", -- 0x1B80
    x"3F",x"3E",x"3E",x"3F",x"3F",x"0F",x"08",x"08", -- 0x1B88
    x"28",x"00",x"08",x"E0",x"C0",x"F0",x"B0",x"B0", -- 0x1B90
    x"F0",x"F0",x"F0",x"F0",x"F0",x"C0",x"80",x"80", -- 0x1B98
    x"A0",x"00",x"FE",x"A0",x"FC",x"FE",x"A0",x"FC", -- 0x1BA0
    x"A0",x"A0",x"FC",x"A0",x"A0",x"E0",x"A0",x"20", -- 0x1BA8
    x"78",x"A0",x"20",x"A0",x"A0",x"20",x"A0",x"A0", -- 0x1BB0
    x"20",x"60",x"A0",x"6A",x"A0",x"A0",x"20",x"A0", -- 0x1BB8
    x"A0",x"A0",x"EC",x"A0",x"A0",x"60",x"A0",x"20", -- 0x1BC0
    x"A0",x"A0",x"20",x"A0",x"A0",x"7C",x"A0",x"A0", -- 0x1BC8
    x"20",x"60",x"FB",x"A0",x"EC",x"FB",x"A0",x"EC", -- 0x1BD0
    x"A0",x"20",x"A0",x"A0",x"20",x"60",x"CC",x"8F", -- 0x1BD8
    x"E8",x"0A",x"50",x"50",x"50",x"50",x"0A",x"0A", -- 0x1BE0
    x"0A",x"0A",x"50",x"50",x"50",x"50",x"00",x"00", -- 0x1BE8
    x"00",x"00",x"50",x"50",x"50",x"50",x"00",x"00", -- 0x1BF0
    x"00",x"00",x"50",x"50",x"50",x"50",x"00",x"00", -- 0x1BF8
    x"00",x"00",x"50",x"50",x"50",x"50",x"08",x"08", -- 0x1C00
    x"02",x"02",x"02",x"02",x"08",x"08",x"50",x"50", -- 0x1C08
    x"50",x"50",x"05",x"05",x"05",x"05",x"20",x"20", -- 0x1C10
    x"80",x"80",x"80",x"80",x"20",x"20",x"05",x"05", -- 0x1C18
    x"05",x"05",x"40",x"40",x"40",x"4A",x"6A",x"6F", -- 0x1C20
    x"6A",x"4A",x"40",x"40",x"40",x"00",x"00",x"00", -- 0x1C28
    x"00",x"00",x"10",x"10",x"10",x"10",x"90",x"90", -- 0x1C30
    x"90",x"10",x"10",x"10",x"10",x"00",x"00",x"00", -- 0x1C38
    x"00",x"00",x"40",x"40",x"40",x"40",x"42",x"4A", -- 0x1C40
    x"6B",x"6F",x"4B",x"4A",x"42",x"40",x"40",x"40", -- 0x1C48
    x"40",x"00",x"01",x"01",x"01",x"01",x"81",x"A1", -- 0x1C50
    x"E9",x"F9",x"E9",x"A1",x"81",x"01",x"01",x"01", -- 0x1C58
    x"01",x"00",x"01",x"05",x"15",x"19",x"5D",x"55", -- 0x1C60
    x"33",x"33",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C68
    x"00",x"00",x"00",x"40",x"50",x"90",x"D4",x"54", -- 0x1C70
    x"30",x"30",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C78
    x"00",x"00",x"01",x"05",x"17",x"5F",x"17",x"05", -- 0x1C80
    x"21",x"80",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C88
    x"00",x"00",x"00",x"40",x"50",x"D4",x"50",x"40", -- 0x1C90
    x"20",x"08",x"30",x"FC",x"B8",x"B8",x"FC",x"EC", -- 0x1C98
    x"EC",x"FC",x"FC",x"88",x"88",x"00",x"00",x"00", -- 0x1CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC0
    x"00",x"00",x"10",x"38",x"54",x"EE",x"7C",x"82", -- 0x1CC8
    x"44",x"00",x"82",x"7C",x"D6",x"FE",x"7C",x"54", -- 0x1CD0
    x"92",x"00",x"00",x"38",x"7C",x"D6",x"EE",x"54", -- 0x1CD8
    x"82",x"00",x"00",x"38",x"7C",x"D6",x"FE",x"44", -- 0x1CE0
    x"28",x"00",x"82",x"7C",x"D6",x"FE",x"7C",x"AA", -- 0x1CE8
    x"54",x"00",x"10",x"38",x"54",x"EE",x"7C",x"44", -- 0x1CF0
    x"82",x"00",x"44",x"44",x"20",x"20",x"44",x"44", -- 0x1CF8
    x"00",x"00",x"44",x"64",x"74",x"64",x"44",x"00", -- 0x1D00
    x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x1D08
    x"F0",x"00",x"38",x"2C",x"FA",x"AF",x"EB",x"AE", -- 0x1D10
    x"38",x"2C",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0", -- 0x1D18
    x"C0",x"C0",x"40",x"08",x"00",x"30",x"03",x"80", -- 0x1D20
    x"04",x"20",x"03",x"10",x"08",x"29",x"C8",x"2C", -- 0x1D28
    x"04",x"40",x"40",x"08",x"00",x"00",x"31",x"00", -- 0x1D30
    x"00",x"00",x"40",x"0C",x"00",x"02",x"80",x"04", -- 0x1D38
    x"00",x"00",x"00",x"30",x"00",x"01",x"00",x"00", -- 0x1D40
    x"08",x"C0",x"00",x"02",x"00",x"10",x"00",x"0C", -- 0x1D48
    x"00",x"80",x"00",x"0C",x"C0",x"00",x"00",x"2E", -- 0x1D50
    x"0A",x"0A",x"0A",x"4A",x"00",x"00",x"01",x"30", -- 0x1D58
    x"00",x"00",x"00",x"40",x"03",x"00",x"00",x"04", -- 0x1D60
    x"80",x"A0",x"80",x"C0",x"00",x"00",x"0C",x"00", -- 0x1D68
    x"00",x"40",x"00",x"00",x"00",x"00",x"00",x"08", -- 0x1D70
    x"0A",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D78
    x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"AA", -- 0x1D80
    x"AA",x"AA",x"02",x"00",x"00",x"00",x"00",x"00", -- 0x1D88
    x"00",x"00",x"00",x"0A",x"2A",x"A9",x"A5",x"95", -- 0x1D90
    x"55",x"95",x"A5",x"A9",x"2A",x"0A",x"00",x"00", -- 0x1D98
    x"00",x"00",x"30",x"AA",x"AA",x"55",x"5F",x"73", -- 0x1DA0
    x"CF",x"7C",x"5F",x"51",x"A2",x"A2",x"01",x"00", -- 0x1DA8
    x"00",x"00",x"C3",x"AA",x"AA",x"55",x"F5",x"3D", -- 0x1DB0
    x"CF",x"FD",x"F5",x"55",x"AA",x"AA",x"54",x"54", -- 0x1DB8
    x"55",x"15",x"0C",x"AA",x"AA",x"5A",x"5A",x"5A", -- 0x1DC0
    x"5A",x"5A",x"5A",x"5A",x"AA",x"AA",x"00",x"00", -- 0x1DC8
    x"00",x"00",x"00",x"00",x"A8",x"00",x"55",x"00", -- 0x1DD0
    x"55",x"00",x"55",x"00",x"A8",x"00",x"00",x"00", -- 0x1DD8
    x"00",x"00",x"15",x"05",x"05",x"15",x"1F",x"15", -- 0x1DE0
    x"00",x"00",x"40",x"40",x"50",x"55",x"FF",x"55", -- 0x1DE8
    x"00",x"00",x"00",x"00",x"00",x"55",x"FF",x"55", -- 0x1DF0
    x"00",x"00",x"00",x"00",x"00",x"55",x"FD",x"55", -- 0x1DF8
    x"00",x"00",x"F0",x"C3",x"C3",x"F3",x"33",x"33", -- 0x1E00
    x"F0",x"00",x"C3",x"0C",x"0C",x"0C",x"0C",x"0C", -- 0x1E08
    x"C3",x"00",x"0F",x"CC",x"CC",x"CF",x"CC",x"CC", -- 0x1E10
    x"0C",x"00",x"0F",x"CC",x"CC",x"0F",x"CC",x"CC", -- 0x1E18
    x"CF",x"00",x"00",x"30",x"30",x"00",x"30",x"30", -- 0x1E20
    x"00",x"00",x"FC",x"CC",x"CC",x"CC",x"CC",x"CC", -- 0x1E28
    x"FC",x"00",x"30",x"F0",x"30",x"30",x"30",x"30", -- 0x1E30
    x"FC",x"00",x"30",x"CC",x"0C",x"0C",x"30",x"C0", -- 0x1E38
    x"FC",x"00",x"FC",x"0C",x"0C",x"30",x"0C",x"CC", -- 0x1E40
    x"30",x"00",x"CC",x"CC",x"CC",x"FC",x"0C",x"0C", -- 0x1E48
    x"0C",x"00",x"FC",x"C0",x"F0",x"0C",x"0C",x"CC", -- 0x1E50
    x"30",x"00",x"30",x"CC",x"C0",x"F0",x"CC",x"CC", -- 0x1E58
    x"30",x"00",x"FC",x"0C",x"0C",x"30",x"30",x"30", -- 0x1E60
    x"30",x"00",x"30",x"CC",x"CC",x"30",x"CC",x"CC", -- 0x1E68
    x"30",x"00",x"30",x"CC",x"CC",x"3C",x"0C",x"0C", -- 0x1E70
    x"0C",x"00",x"30",x"30",x"30",x"FC",x"FC",x"FC", -- 0x1E78
    x"FC",x"CC",x"F0",x"F0",x"F0",x"F0",x"00",x"00", -- 0x1E80
    x"00",x"00",x"40",x"00",x"00",x"00",x"00",x"00", -- 0x1E88
    x"00",x"00",x"80",x"01",x"00",x"01",x"8C",x"00", -- 0x1E90
    x"DC",x"E6",x"F0",x"FA",x"F9",x"F8",x"F7",x"F6", -- 0x1E98
    x"F5",x"F4",x"F3",x"F2",x"F1",x"F0",x"EF",x"EE", -- 0x1EA0
    x"ED",x"EC",x"EB",x"EA",x"E9",x"E8",x"E7",x"E6", -- 0x1EA8
    x"00",x"AA",x"AF",x"B4",x"BE",x"C8",x"D2",x"D7", -- 0x1EB0
    x"DC",x"E1",x"E6",x"EB",x"F0",x"F5",x"FA",x"FF", -- 0x1EB8
    x"00",x"FF",x"FA",x"F5",x"F0",x"EB",x"E6",x"E1", -- 0x1EC0
    x"DC",x"D7",x"D2",x"C8",x"BE",x"B4",x"AF",x"AA", -- 0x1EC8
    x"00",x"F0",x"01",x"DC",x"01",x"E6",x"01",x"D2", -- 0x1ED0
    x"01",x"E1",x"01",x"D7",x"01",x"E6",x"01",x"D2", -- 0x1ED8
    x"01",x"00",x"DC",x"D7",x"D6",x"D4",x"D2",x"D0", -- 0x1EE0
    x"CE",x"CC",x"CA",x"C8",x"C6",x"C3",x"C0",x"BE", -- 0x1EE8
    x"BC",x"B9",x"B6",x"B4",x"AF",x"AA",x"A5",x"A0", -- 0x1EF0
    x"00",x"BE",x"C3",x"C8",x"CD",x"D2",x"D7",x"DC", -- 0x1EF8
    x"E1",x"E6",x"F0",x"F5",x"FA",x"00",x"80",x"00", -- 0x1F00
    x"B4",x"B2",x"B0",x"AE",x"AC",x"AA",x"AC",x"AE", -- 0x1F08
    x"B0",x"B2",x"00",x"01",x"CD",x"01",x"C8",x"01", -- 0x1F10
    x"C3",x"01",x"BE",x"01",x"B4",x"01",x"8C",x"01", -- 0x1F18
    x"00",x"01",x"01",x"00",x"3C",x"01",x"00",x"01", -- 0x1F20
    x"02",x"02",x"02",x"02",x"02",x"02",x"03",x"03", -- 0x1F28
    x"03",x"03",x"04",x"04",x"04",x"04",x"04",x"03", -- 0x1F30
    x"03",x"03",x"03",x"02",x"02",x"01",x"01",x"00", -- 0x1F38
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x1F40
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00", -- 0x1F48
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x1F50
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00", -- 0x1F58
    x"01",x"02",x"01",x"02",x"01",x"02",x"01",x"02", -- 0x1F60
    x"01",x"02",x"01",x"02",x"01",x"02",x"01",x"01", -- 0x1F68
    x"00",x"03",x"03",x"03",x"03",x"03",x"03",x"03", -- 0x1F70
    x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03", -- 0x1F78
    x"03",x"03",x"03",x"03",x"03",x"03",x"01",x"00", -- 0x1F80
    x"04",x"04",x"04",x"04",x"03",x"03",x"03",x"03", -- 0x1F88
    x"03",x"03",x"03",x"01",x"00",x"01",x"00",x"03", -- 0x1F90
    x"03",x"03",x"04",x"04",x"04",x"03",x"03",x"03", -- 0x1F98
    x"01",x"00",x"01",x"0F",x"01",x"0F",x"01",x"0F", -- 0x1FA0
    x"01",x"0F",x"01",x"0F",x"01",x"0F",x"01",x"00", -- 0x1FA8
    x"02",x"19",x"00",x"02",x"09",x"0C",x"0C",x"20", -- 0x1FB0
    x"08",x"09",x"0E",x"04",x"0F",x"12",x"06",x"06", -- 0x1FB8
    x"00",x"01",x"0E",x"04",x"19",x"20",x"06",x"09", -- 0x1FC0
    x"0E",x"0B",x"05",x"0C",x"00",x"0A",x"05",x"06", -- 0x1FC8
    x"06",x"20",x"02",x"12",x"15",x"05",x"14",x"14", -- 0x1FD0
    x"05",x"00",x"05",x"12",x"09",x"03",x"20",x"03", -- 0x1FD8
    x"0F",x"14",x"14",x"0F",x"0E",x"00",x"0D",x"01", -- 0x1FE0
    x"12",x"0B",x"20",x"13",x"03",x"0F",x"14",x"14", -- 0x1FE8
    x"00",x"0A",x"09",x"0D",x"0D",x"19",x"20",x"13", -- 0x1FF0
    x"0E",x"19",x"04",x"05",x"12",x"00",x"FF",x"AA"  -- 0x1FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
