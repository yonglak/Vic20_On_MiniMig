-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity cart_rom is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of cart_rom is


  type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"11",x"A0",x"11",x"A0",x"41",x"30",x"C3",x"C2", -- 0x0000 --41
    x"CD",x"02",x"BB",x"5A",x"30",x"5F",x"EE",x"3D", -- 0x0008
    x"A8",x"20",x"52",x"FD",x"20",x"F9",x"FD",x"20", -- 0x0010
    x"18",x"E5",x"78",x"D8",x"20",x"68",x"AE",x"CA", -- 0x0018
    x"9A",x"A9",x"8C",x"8D",x"05",x"90",x"A9",x"96", -- 0x0020
    x"8D",x"02",x"90",x"A9",x"7F",x"8D",x"1E",x"91", -- 0x0028
    x"A9",x"17",x"8D",x"03",x"90",x"E8",x"8A",x"95", -- 0x0030
    x"00",x"CA",x"D0",x"FB",x"A9",x"00",x"8D",x"05", -- 0x0038
    x"01",x"8D",x"04",x"01",x"A0",x"ED",x"A9",x"00", -- 0x0040
    x"99",x"00",x"00",x"88",x"D0",x"FA",x"A9",x"00", -- 0x0048
    x"85",x"00",x"A8",x"A2",x"16",x"99",x"00",x"02", -- 0x0050
    x"C8",x"18",x"69",x"0B",x"CA",x"D0",x"F6",x"E6", -- 0x0058
    x"00",x"A5",x"00",x"C9",x"0B",x"D0",x"EC",x"A9", -- 0x0060
    x"FF",x"A2",x"16",x"99",x"00",x"02",x"99",x"08", -- 0x0068
    x"02",x"C8",x"F0",x"03",x"CA",x"10",x"F4",x"A9", -- 0x0070
    x"96",x"A0",x"00",x"84",x"FB",x"85",x"FC",x"99", -- 0x0078
    x"DA",x"03",x"A5",x"FB",x"99",x"BC",x"03",x"18", -- 0x0080
    x"69",x"16",x"85",x"FB",x"A5",x"FC",x"69",x"00", -- 0x0088
    x"C8",x"C0",x"1A",x"D0",x"E8",x"A9",x"00",x"85", -- 0x0090
    x"F7",x"A9",x"10",x"A0",x"00",x"85",x"F8",x"99", -- 0x0098
    x"9E",x"03",x"A5",x"F7",x"99",x"80",x"03",x"18", -- 0x00A0
    x"69",x"B0",x"85",x"F7",x"A5",x"F8",x"69",x"00", -- 0x00A8
    x"C8",x"C0",x"18",x"D0",x"E8",x"A9",x"80",x"85", -- 0x00B0
    x"F7",x"A9",x"9E",x"85",x"F9",x"A9",x"03",x"85", -- 0x00B8
    x"F8",x"85",x"FA",x"A9",x"BC",x"85",x"FB",x"A9", -- 0x00C0
    x"DA",x"85",x"FD",x"A9",x"03",x"85",x"FC",x"85", -- 0x00C8
    x"FE",x"A9",x"0E",x"8D",x"0F",x"90",x"A9",x"2F", -- 0x00D0
    x"8D",x"0E",x"90",x"A9",x"01",x"8D",x"02",x"01", -- 0x00D8
    x"20",x"9D",x"A7",x"A0",x"07",x"A9",x"00",x"99", -- 0x00E0
    x"EC",x"00",x"88",x"10",x"FA",x"A2",x"1D",x"BD", -- 0x00E8
    x"2C",x"B0",x"9D",x"E1",x"1F",x"CA",x"10",x"F7", -- 0x00F0
    x"A2",x"1D",x"BD",x"0E",x"B0",x"95",x"AB",x"BD", -- 0x00F8
    x"2C",x"B0",x"95",x"C9",x"CA",x"10",x"F3",x"A9", -- 0x0100
    x"0F",x"A2",x"00",x"A0",x"16",x"20",x"4F",x"AE", -- 0x0108
    x"A2",x"00",x"A0",x"00",x"A9",x"07",x"20",x"4F", -- 0x0110
    x"AE",x"A2",x"0A",x"A0",x"0A",x"20",x"4F",x"AE", -- 0x0118
    x"A0",x"C8",x"A9",x"00",x"99",x"00",x"00",x"88", -- 0x0120
    x"D0",x"FA",x"A2",x"1D",x"B5",x"C9",x"F0",x"0A", -- 0x0128
    x"BD",x"0E",x"B0",x"95",x"AB",x"BD",x"2C",x"B0", -- 0x0130
    x"95",x"C9",x"CA",x"10",x"EF",x"A9",x"01",x"85", -- 0x0138
    x"1E",x"A9",x"23",x"85",x"1F",x"A2",x"28",x"86", -- 0x0140
    x"25",x"A2",x"1D",x"86",x"20",x"20",x"68",x"AE", -- 0x0148
    x"20",x"4F",x"AD",x"20",x"D1",x"AB",x"20",x"48", -- 0x0150
    x"AC",x"20",x"B5",x"A9",x"20",x"F5",x"A5",x"20", -- 0x0158
    x"7C",x"A6",x"20",x"8E",x"A4",x"20",x"C9",x"A4", -- 0x0160
    x"20",x"77",x"A1",x"20",x"D3",x"A5",x"20",x"FA", -- 0x0168
    x"A4",x"20",x"A1",x"AC",x"4C",x"5C",x"A1",x"C6", -- 0x0170
    x"27",x"10",x"40",x"A9",x"05",x"85",x"27",x"20", -- 0x0178
    x"3A",x"A2",x"20",x"20",x"A7",x"A2",x"02",x"86", -- 0x0180
    x"21",x"A6",x"20",x"B5",x"C9",x"F0",x"2D",x"95", -- 0x0188
    x"C9",x"85",x"0E",x"B5",x"6E",x"D0",x"06",x"20", -- 0x0190
    x"C2",x"A1",x"20",x"E1",x"A1",x"A6",x"20",x"CA", -- 0x0198
    x"10",x"13",x"A2",x"1D",x"C6",x"1F",x"D0",x"0D", -- 0x01A0
    x"A5",x"1E",x"49",x"FF",x"18",x"69",x"01",x"85", -- 0x01A8
    x"1E",x"A9",x"23",x"85",x"1F",x"86",x"20",x"C6", -- 0x01B0
    x"21",x"10",x"D0",x"60",x"20",x"98",x"A7",x"4C", -- 0x01B8
    x"9D",x"A1",x"BD",x"0E",x"B0",x"85",x"00",x"A4", -- 0x01C0
    x"1E",x"10",x"09",x"18",x"65",x"1F",x"38",x"E9", -- 0x01C8
    x"01",x"4C",x"DC",x"A1",x"A9",x"23",x"38",x"E5", -- 0x01D0
    x"1F",x"18",x"65",x"00",x"95",x"AB",x"85",x"0D", -- 0x01D8
    x"60",x"29",x"01",x"18",x"7D",x"D2",x"AF",x"4C", -- 0x01E0
    x"C6",x"AE",x"A6",x"96",x"20",x"C2",x"A1",x"B5", -- 0x01E8
    x"C9",x"18",x"69",x"01",x"95",x"C9",x"85",x"0E", -- 0x01F0
    x"DD",x"2C",x"B0",x"F0",x"0C",x"20",x"E1",x"A1", -- 0x01F8
    x"4C",x"E9",x"A2",x"20",x"98",x"A7",x"4C",x"E9", -- 0x0200
    x"A2",x"A6",x"96",x"A9",x"00",x"95",x"6E",x"A4", -- 0x0208
    x"95",x"99",x"8C",x"00",x"10",x"E7",x"20",x"B0", -- 0x0210
    x"AE",x"A6",x"96",x"B4",x"C9",x"B5",x"AB",x"AA", -- 0x0218
    x"A9",x"0A",x"20",x"C2",x"AE",x"A6",x"95",x"B5", -- 0x0220
    x"8C",x"09",x"E0",x"95",x"8C",x"A4",x"96",x"99", -- 0x0228
    x"6E",x"00",x"A9",x"0F",x"99",x"C9",x"00",x"4C", -- 0x0230
    x"EA",x"A1",x"A9",x"00",x"85",x"A3",x"A2",x"08", -- 0x0238
    x"86",x"95",x"B5",x"8C",x"F0",x"BD",x"29",x"1F", -- 0x0240
    x"85",x"96",x"B5",x"8C",x"29",x"E0",x"C9",x"E0", -- 0x0248
    x"F0",x"E5",x"20",x"C8",x"A6",x"A6",x"95",x"A4", -- 0x0250
    x"96",x"B9",x"6E",x"00",x"29",x"7F",x"38",x"E9", -- 0x0258
    x"01",x"D0",x"03",x"4C",x"09",x"A3",x"85",x"99", -- 0x0260
    x"B9",x"6E",x"00",x"29",x"80",x"85",x"98",x"05", -- 0x0268
    x"99",x"99",x"6E",x"00",x"B5",x"8C",x"4A",x"4A", -- 0x0270
    x"4A",x"4A",x"4A",x"38",x"E9",x"01",x"0A",x"AA", -- 0x0278
    x"BD",x"8E",x"B0",x"85",x"02",x"BD",x"98",x"B0", -- 0x0280
    x"85",x"04",x"E8",x"BD",x"8E",x"B0",x"85",x"03", -- 0x0288
    x"BD",x"98",x"B0",x"85",x"05",x"A6",x"96",x"A4", -- 0x0290
    x"99",x"B5",x"C9",x"18",x"71",x"04",x"C9",x"96", -- 0x0298
    x"90",x"03",x"4C",x"16",x"A2",x"95",x"C9",x"85", -- 0x02A0
    x"0E",x"4A",x"C5",x"A3",x"90",x"02",x"85",x"A3", -- 0x02A8
    x"A5",x"98",x"30",x"07",x"B1",x"02",x"F0",x"05", -- 0x02B0
    x"A9",x"FF",x"2C",x"B1",x"02",x"85",x"00",x"B5", -- 0x02B8
    x"AB",x"18",x"65",x"00",x"C9",x"54",x"90",x"03", -- 0x02C0
    x"4C",x"16",x"A2",x"95",x"AB",x"85",x"0D",x"86", -- 0x02C8
    x"21",x"20",x"E1",x"A1",x"A6",x"21",x"B5",x"C9", -- 0x02D0
    x"C9",x"91",x"90",x"0D",x"B5",x"AB",x"38",x"E5", -- 0x02D8
    x"25",x"C9",x"FD",x"B0",x"15",x"C9",x"05",x"90", -- 0x02E0
    x"11",x"A6",x"95",x"CA",x"30",x"03",x"4C",x"40", -- 0x02E8
    x"A2",x"A9",x"00",x"38",x"E5",x"A3",x"8D",x"0A", -- 0x02F0
    x"90",x"60",x"A5",x"9C",x"D0",x"07",x"A9",x"0B", -- 0x02F8
    x"85",x"9C",x"20",x"DD",x"A3",x"4C",x"E9",x"A2", -- 0x0300
    x"60",x"C0",x"10",x"B0",x"1C",x"A5",x"A4",x"C9", -- 0x0308
    x"04",x"90",x"23",x"A2",x"01",x"20",x"FF",x"AD", -- 0x0310
    x"F0",x"F3",x"48",x"A2",x"07",x"20",x"FF",x"AD", -- 0x0318
    x"29",x"80",x"85",x"01",x"68",x"AA",x"4C",x"50", -- 0x0320
    x"A3",x"C0",x"10",x"90",x"09",x"C0",x"16",x"B0", -- 0x0328
    x"05",x"A2",x"04",x"4C",x"50",x"A3",x"B9",x"AB", -- 0x0330
    x"00",x"38",x"E5",x"25",x"A2",x"01",x"C9",x"14", -- 0x0338
    x"90",x"0E",x"C9",x"EB",x"B0",x"0A",x"E8",x"C9", -- 0x0340
    x"1E",x"90",x"05",x"C9",x"E1",x"B0",x"01",x"E8", -- 0x0348
    x"86",x"00",x"E8",x"8A",x"0A",x"0A",x"0A",x"0A", -- 0x0350
    x"0A",x"85",x"21",x"05",x"96",x"A6",x"95",x"95", -- 0x0358
    x"8C",x"A6",x"00",x"BD",x"89",x"B0",x"A6",x"A4", -- 0x0360
    x"E0",x"04",x"90",x"0B",x"A6",x"96",x"E0",x"10", -- 0x0368
    x"B0",x"05",x"05",x"01",x"4C",x"81",x"A3",x"A6", -- 0x0370
    x"96",x"B4",x"AB",x"C4",x"25",x"B0",x"02",x"09", -- 0x0378
    x"80",x"95",x"6E",x"85",x"01",x"A5",x"95",x"C9", -- 0x0380
    x"08",x"F0",x"05",x"A6",x"95",x"4C",x"57",x"A2", -- 0x0388
    x"A2",x"07",x"B5",x"8C",x"F0",x"03",x"20",x"A4", -- 0x0390
    x"A3",x"CA",x"B5",x"8C",x"F0",x"ED",x"20",x"A4", -- 0x0398
    x"A3",x"4C",x"8B",x"A3",x"29",x"E0",x"C9",x"E0", -- 0x03A0
    x"F0",x"12",x"B5",x"8C",x"29",x"1F",x"A8",x"A5", -- 0x03A8
    x"01",x"99",x"6E",x"00",x"B5",x"8C",x"29",x"1F", -- 0x03B0
    x"05",x"21",x"95",x"8C",x"60",x"A5",x"2B",x"F0", -- 0x03B8
    x"FB",x"A2",x"1D",x"86",x"21",x"B5",x"C9",x"F0", -- 0x03C0
    x"76",x"38",x"E5",x"2A",x"C9",x"03",x"90",x"04", -- 0x03C8
    x"C9",x"FA",x"90",x"6B",x"B5",x"AB",x"38",x"E5", -- 0x03D0
    x"29",x"C9",x"FC",x"90",x"62",x"20",x"B0",x"AE", -- 0x03D8
    x"A0",x"08",x"B9",x"8C",x"00",x"F0",x"06",x"29", -- 0x03E0
    x"1F",x"C5",x"21",x"F0",x"05",x"88",x"10",x"F2", -- 0x03E8
    x"30",x"13",x"A9",x"00",x"99",x"8C",x"00",x"95", -- 0x03F0
    x"6E",x"C0",x"06",x"B0",x"4B",x"BD",x"F0",x"AF", -- 0x03F8
    x"A2",x"00",x"20",x"F7",x"AC",x"A6",x"21",x"B4", -- 0x0400
    x"C9",x"A9",x"00",x"95",x"C9",x"95",x"6E",x"B5", -- 0x0408
    x"AB",x"AA",x"A9",x"0A",x"20",x"C2",x"AE",x"A2", -- 0x0410
    x"07",x"B5",x"53",x"F0",x"06",x"CA",x"10",x"F9", -- 0x0418
    x"4C",x"F8",x"A0",x"A5",x"0D",x"95",x"5B",x"A5", -- 0x0420
    x"0E",x"95",x"63",x"A9",x"03",x"95",x"53",x"A6", -- 0x0428
    x"21",x"BD",x"F0",x"AF",x"A2",x"00",x"20",x"F7", -- 0x0430
    x"AC",x"20",x"C9",x"A4",x"4C",x"B8",x"A6",x"A6", -- 0x0438
    x"21",x"CA",x"30",x"03",x"4C",x"C3",x"A3",x"60", -- 0x0440
    x"E6",x"9A",x"C0",x"08",x"D0",x"AF",x"A9",x"FF", -- 0x0448
    x"85",x"A5",x"A9",x"03",x"85",x"A6",x"A4",x"9A", -- 0x0450
    x"BE",x"BA",x"AF",x"86",x"05",x"B9",x"C2",x"AF", -- 0x0458
    x"85",x"04",x"20",x"F7",x"AC",x"A2",x"1C",x"A0", -- 0x0460
    x"A8",x"A9",x"04",x"85",x"22",x"A9",x"00",x"85", -- 0x0468
    x"23",x"A9",x"FF",x"85",x"9B",x"F8",x"A5",x"04", -- 0x0470
    x"18",x"69",x"60",x"85",x"04",x"A5",x"05",x"69", -- 0x0478
    x"00",x"85",x"05",x"D8",x"A9",x"01",x"20",x"80", -- 0x0480
    x"AD",x"A6",x"21",x"4C",x"05",x"A4",x"C6",x"6B", -- 0x0488
    x"10",x"B5",x"A9",x"0A",x"85",x"6B",x"A2",x"07", -- 0x0490
    x"86",x"21",x"B5",x"53",x"F0",x"25",x"B5",x"63", -- 0x0498
    x"85",x"0E",x"B5",x"5B",x"85",x"0D",x"A9",x"0B", -- 0x04A0
    x"38",x"F5",x"53",x"20",x"C6",x"AE",x"A6",x"21", -- 0x04A8
    x"B5",x"53",x"0A",x"0A",x"0A",x"0A",x"18",x"69", -- 0x04B0
    x"7F",x"8D",x"0D",x"90",x"D6",x"53",x"D0",x"03", -- 0x04B8
    x"20",x"AA",x"AE",x"A6",x"21",x"CA",x"10",x"D0", -- 0x04C0
    x"60",x"A9",x"00",x"85",x"A4",x"A2",x"1D",x"B5", -- 0x04C8
    x"C9",x"F0",x"02",x"E6",x"A4",x"CA",x"10",x"F7", -- 0x04D0
    x"A5",x"A4",x"C9",x"06",x"B0",x"04",x"A9",x"01", -- 0x04D8
    x"85",x"A7",x"A5",x"A4",x"D0",x"E2",x"A5",x"9C", -- 0x04E0
    x"F0",x"01",x"60",x"A6",x"25",x"A0",x"98",x"A9", -- 0x04E8
    x"0A",x"20",x"C2",x"AE",x"20",x"B8",x"A6",x"4C", -- 0x04F0
    x"29",x"AC",x"C6",x"A5",x"D0",x"CA",x"C6",x"A6", -- 0x04F8
    x"10",x"C6",x"A9",x"01",x"85",x"A5",x"A9",x"00", -- 0x0500
    x"85",x"A6",x"A5",x"A7",x"D0",x"0C",x"A6",x"E7", -- 0x0508
    x"B4",x"6C",x"BE",x"77",x"B0",x"20",x"FF",x"AD", -- 0x0510
    x"D0",x"AE",x"A6",x"E7",x"B5",x"EA",x"C9",x"06", -- 0x0518
    x"90",x"03",x"A2",x"00",x"2C",x"A2",x"01",x"20", -- 0x0520
    x"FF",x"AD",x"D0",x"10",x"A9",x"1C",x"85",x"00", -- 0x0528
    x"A5",x"E6",x"05",x"E5",x"F0",x"0A",x"A0",x"01", -- 0x0530
    x"B5",x"8C",x"F0",x"39",x"A9",x"16",x"85",x"00", -- 0x0538
    x"A2",x"05",x"B5",x"8C",x"F0",x"04",x"CA",x"10", -- 0x0540
    x"F9",x"60",x"86",x"95",x"A2",x"1B",x"BC",x"4A", -- 0x0548
    x"B0",x"C4",x"00",x"B0",x"0A",x"B9",x"C9",x"00", -- 0x0550
    x"F0",x"05",x"B9",x"6E",x"00",x"F0",x"04",x"CA", -- 0x0558
    x"10",x"EC",x"60",x"84",x"96",x"98",x"09",x"20", -- 0x0560
    x"A6",x"95",x"95",x"8C",x"A9",x"12",x"19",x"A2", -- 0x0568
    x"B0",x"99",x"6E",x"00",x"60",x"A2",x"00",x"20", -- 0x0570
    x"FF",x"AD",x"18",x"69",x"1C",x"A8",x"A2",x"08", -- 0x0578
    x"B9",x"C9",x"00",x"F0",x"B7",x"B5",x"8C",x"D0", -- 0x0580
    x"B3",x"A9",x"01",x"85",x"9A",x"86",x"95",x"84", -- 0x0588
    x"96",x"20",x"63",x"A5",x"A5",x"96",x"38",x"E9", -- 0x0590
    x"1C",x"AA",x"A0",x"07",x"84",x"95",x"0A",x"0A", -- 0x0598
    x"09",x"03",x"85",x"00",x"A9",x"02",x"85",x"01", -- 0x05A0
    x"A6",x"00",x"BC",x"CA",x"AF",x"F0",x"C5",x"B9", -- 0x05A8
    x"C9",x"00",x"F0",x"17",x"B9",x"6E",x"00",x"D0", -- 0x05B0
    x"12",x"A6",x"95",x"B5",x"8C",x"D0",x"0C",x"20", -- 0x05B8
    x"63",x"A5",x"A5",x"9A",x"0A",x"85",x"9A",x"C6", -- 0x05C0
    x"95",x"C6",x"01",x"A5",x"01",x"F0",x"A5",x"C6", -- 0x05C8
    x"00",x"10",x"D5",x"A5",x"9B",x"F0",x"9D",x"C6", -- 0x05D0
    x"9B",x"D0",x"99",x"A2",x"28",x"86",x"0D",x"A0", -- 0x05D8
    x"A8",x"84",x"0E",x"A9",x"16",x"20",x"C6",x"AE", -- 0x05E0
    x"A5",x"0D",x"38",x"E9",x"04",x"C9",x"18",x"F0", -- 0x05E8
    x"83",x"85",x"0D",x"10",x"EE",x"A5",x"9C",x"D0", -- 0x05F0
    x"57",x"C6",x"26",x"10",x"52",x"A9",x"05",x"85", -- 0x05F8
    x"26",x"20",x"22",x"AE",x"A5",x"25",x"A6",x"0A", -- 0x0600
    x"F0",x"0B",x"A6",x"08",x"D0",x"10",x"38",x"E9", -- 0x0608
    x"01",x"10",x"09",x"30",x"09",x"18",x"69",x"01", -- 0x0610
    x"C9",x"52",x"F0",x"02",x"85",x"25",x"A5",x"2B", -- 0x0618
    x"D0",x"1D",x"A5",x"0C",x"F0",x"06",x"A9",x"00", -- 0x0620
    x"85",x"6D",x"F0",x"13",x"A5",x"6D",x"D0",x"0F", -- 0x0628
    x"E6",x"6D",x"A5",x"25",x"18",x"69",x"03",x"85", -- 0x0630
    x"29",x"85",x"2B",x"A9",x"98",x"85",x"2A",x"A0", -- 0x0638
    x"98",x"A6",x"25",x"A5",x"2B",x"F0",x"03",x"A9", -- 0x0640
    x"11",x"2C",x"A9",x"10",x"4C",x"C2",x"AE",x"60", -- 0x0648
    x"C6",x"9D",x"10",x"FB",x"A9",x"0F",x"85",x"9D", -- 0x0650
    x"A2",x"07",x"20",x"FF",x"AD",x"8D",x"0D",x"90", -- 0x0658
    x"20",x"FF",x"AD",x"8D",x"0A",x"90",x"CE",x"0E", -- 0x0660
    x"90",x"A6",x"9C",x"BD",x"AE",x"AF",x"A6",x"25", -- 0x0668
    x"A0",x"98",x"20",x"C2",x"AE",x"C6",x"9C",x"D0", -- 0x0670
    x"D6",x"4C",x"11",x"AA",x"20",x"8B",x"A6",x"20", -- 0x0678
    x"8B",x"A6",x"20",x"8B",x"A6",x"20",x"8B",x"A6", -- 0x0680
    x"4C",x"BD",x"A3",x"A5",x"2B",x"F0",x"C0",x"C6", -- 0x0688
    x"28",x"10",x"BC",x"A9",x"01",x"85",x"28",x"A5", -- 0x0690
    x"2A",x"4A",x"18",x"69",x"AF",x"8D",x"0B",x"90", -- 0x0698
    x"A5",x"29",x"85",x"0D",x"A5",x"2A",x"85",x"0E", -- 0x06A0
    x"38",x"E9",x"01",x"C9",x"0F",x"F0",x"09",x"85", -- 0x06A8
    x"2A",x"85",x"0E",x"A9",x"12",x"4C",x"C6",x"AE", -- 0x06B0
    x"20",x"B6",x"AE",x"85",x"2B",x"A6",x"29",x"A4", -- 0x06B8
    x"2A",x"F0",x"8C",x"A9",x"13",x"4C",x"C2",x"AE", -- 0x06C0
    x"A6",x"E7",x"B4",x"6C",x"BE",x"77",x"B0",x"CA", -- 0x06C8
    x"20",x"FF",x"AD",x"D0",x"0E",x"A6",x"E7",x"B4", -- 0x06D0
    x"6C",x"BE",x"80",x"B0",x"B5",x"47",x"F0",x"04", -- 0x06D8
    x"CA",x"10",x"F9",x"60",x"86",x"2E",x"A4",x"96", -- 0x06E0
    x"B9",x"C9",x"00",x"F0",x"F6",x"C9",x"7C",x"B0", -- 0x06E8
    x"F2",x"18",x"69",x"0C",x"95",x"3B",x"85",x"0E", -- 0x06F0
    x"B9",x"AB",x"00",x"18",x"69",x"03",x"C9",x"54", -- 0x06F8
    x"B0",x"E1",x"95",x"2F",x"85",x"0D",x"A6",x"96", -- 0x0700
    x"A0",x"01",x"B5",x"AB",x"C5",x"25",x"90",x"07", -- 0x0708
    x"98",x"49",x"FF",x"18",x"69",x"01",x"A8",x"A6", -- 0x0710
    x"2E",x"94",x"47",x"A9",x"14",x"4C",x"C6",x"AE", -- 0x0718
    x"C6",x"A8",x"10",x"BF",x"A9",x"01",x"85",x"A8", -- 0x0720
    x"A6",x"E7",x"B4",x"6C",x"BE",x"80",x"B0",x"86", -- 0x0728
    x"2E",x"B5",x"47",x"F0",x"47",x"B5",x"3B",x"85", -- 0x0730
    x"0E",x"B5",x"2F",x"85",x"0D",x"A9",x"13",x"20", -- 0x0738
    x"C6",x"AE",x"A6",x"2E",x"B5",x"2F",x"30",x"47", -- 0x0740
    x"C9",x"54",x"B0",x"43",x"85",x"0D",x"B5",x"3B", -- 0x0748
    x"18",x"69",x"05",x"C9",x"9C",x"B0",x"38",x"95", -- 0x0750
    x"3B",x"85",x"0E",x"4A",x"85",x"00",x"A9",x"C8", -- 0x0758
    x"38",x"E5",x"00",x"8D",x"0C",x"90",x"A9",x"14", -- 0x0760
    x"20",x"C6",x"AE",x"A6",x"2E",x"B5",x"3B",x"C9", -- 0x0768
    x"93",x"90",x"09",x"B5",x"2F",x"38",x"E5",x"25", -- 0x0770
    x"C9",x"05",x"90",x"06",x"A6",x"2E",x"CA",x"10", -- 0x0778
    x"AE",x"60",x"A9",x"13",x"20",x"C6",x"AE",x"A5", -- 0x0780
    x"9C",x"D0",x"04",x"A9",x"06",x"85",x"9C",x"A6", -- 0x0788
    x"2E",x"20",x"BC",x"AE",x"95",x"47",x"F0",x"E4", -- 0x0790
    x"A9",x"10",x"4C",x"95",x"AE",x"20",x"59",x"AB", -- 0x0798
    x"20",x"68",x"AE",x"20",x"A1",x"AE",x"8D",x"02", -- 0x07A0
    x"01",x"20",x"CC",x"A9",x"A2",x"08",x"A0",x"08", -- 0x07A8
    x"20",x"CD",x"AD",x"31",x"22",x"31",x"2A",x"20", -- 0x07B0
    x"24",x"2D",x"1B",x"22",x"16",x"28",x"2A",x"2E", -- 0x07B8
    x"24",x"2E",x"29",x"22",x"24",x"00",x"A2",x"1C", -- 0x07C0
    x"A0",x"18",x"20",x"CD",x"AD",x"32",x"31",x"27", -- 0x07C8
    x"31",x"1C",x"20",x"31",x"29",x"00",x"A2",x"18", -- 0x07D0
    x"A0",x"30",x"20",x"CD",x"AD",x"28",x"2A",x"2E", -- 0x07D8
    x"24",x"24",x"16",x"1B",x"34",x"00",x"A2",x"14", -- 0x07E0
    x"A0",x"38",x"20",x"CD",x"AD",x"1B",x"2D",x"2A", -- 0x07E8
    x"16",x"2D",x"28",x"22",x"20",x"2D",x"29",x"24", -- 0x07F0
    x"00",x"A2",x"04",x"A0",x"08",x"A9",x"0F",x"20", -- 0x07F8
    x"4F",x"AE",x"A2",x"1D",x"86",x"20",x"BD",x"2C", -- 0x0800
    x"B0",x"18",x"69",x"3C",x"95",x"C9",x"BD",x"0E", -- 0x0808
    x"B0",x"95",x"AB",x"CA",x"10",x"F0",x"A9",x"15", -- 0x0810
    x"85",x"1F",x"A9",x"01",x"85",x"1E",x"20",x"85", -- 0x0818
    x"A1",x"A5",x"20",x"C9",x"1D",x"D0",x"F7",x"A2", -- 0x0820
    x"14",x"A0",x"A0",x"20",x"CD",x"AD",x"23",x"34", -- 0x0828
    x"3C",x"3B",x"36",x"16",x"31",x"22",x"31",x"2A", -- 0x0830
    x"20",x"00",x"A2",x"04",x"A0",x"A8",x"20",x"CD", -- 0x0838
    x"AD",x"31",x"27",x"27",x"16",x"2A",x"20",x"32", -- 0x0840
    x"1E",x"22",x"24",x"16",x"2A",x"2E",x"24",x"2E", -- 0x0848
    x"2A",x"2C",x"2E",x"21",x"16",x"16",x"00",x"A9", -- 0x0850
    x"01",x"8D",x"02",x"01",x"20",x"70",x"AB",x"20", -- 0x0858
    x"E5",x"A9",x"D0",x"0D",x"20",x"22",x"AE",x"A5", -- 0x0860
    x"0C",x"D0",x"F1",x"20",x"59",x"AB",x"4C",x"90", -- 0x0868
    x"A9",x"20",x"A1",x"AE",x"20",x"59",x"AB",x"20", -- 0x0870
    x"08",x"AA",x"20",x"68",x"AE",x"20",x"CC",x"A9", -- 0x0878
    x"A9",x"00",x"8D",x"02",x"01",x"20",x"4F",x"AD", -- 0x0880
    x"A2",x"10",x"A0",x"28",x"20",x"CD",x"AD",x"1B", -- 0x0888
    x"34",x"26",x"24",x"22",x"31",x"2A",x"22",x"16", -- 0x0890
    x"32",x"31",x"30",x"2E",x"00",x"A2",x"10",x"A0", -- 0x0898
    x"38",x"20",x"CD",x"AD",x"1B",x"36",x"26",x"16", -- 0x08A0
    x"16",x"28",x"27",x"31",x"19",x"2E",x"2A",x"00", -- 0x08A8
    x"AD",x"05",x"01",x"85",x"E7",x"18",x"69",x"34", -- 0x08B0
    x"A2",x"1C",x"A0",x"38",x"20",x"C2",x"AE",x"A2", -- 0x08B8
    x"10",x"A0",x"48",x"20",x"CD",x"AD",x"1B",x"38", -- 0x08C0
    x"26",x"27",x"2E",x"2C",x"2E",x"27",x"00",x"AD", -- 0x08C8
    x"04",x"01",x"85",x"EA",x"85",x"EB",x"18",x"69", -- 0x08D0
    x"34",x"A2",x"34",x"A0",x"48",x"20",x"C2",x"AE", -- 0x08D8
    x"A2",x"10",x"A0",x"70",x"20",x"CD",x"AD",x"06", -- 0x08E0
    x"16",x"16",x"16",x"16",x"16",x"04",x"16",x"16", -- 0x08E8
    x"16",x"02",x"16",x"16",x"16",x"01",x"00",x"A2", -- 0x08F0
    x"10",x"A0",x"80",x"20",x"CD",x"AD",x"39",x"33", -- 0x08F8
    x"16",x"16",x"16",x"16",x"38",x"33",x"16",x"16", -- 0x0900
    x"37",x"33",x"16",x"16",x"36",x"33",x"00",x"A2", -- 0x0908
    x"04",x"A0",x"90",x"20",x"CD",x"AD",x"34",x"38", -- 0x0910
    x"33",x"26",x"3B",x"33",x"33",x"16",x"34",x"33", -- 0x0918
    x"33",x"16",x"16",x"3B",x"33",x"16",x"16",x"39", -- 0x0920
    x"33",x"00",x"A9",x"01",x"8D",x"02",x"01",x"20", -- 0x0928
    x"70",x"AB",x"20",x"22",x"AE",x"A5",x"0C",x"F0", -- 0x0930
    x"57",x"20",x"F0",x"A9",x"A6",x"A1",x"85",x"A1", -- 0x0938
    x"E0",x"01",x"F0",x"1F",x"C9",x"00",x"F0",x"1B", -- 0x0940
    x"A5",x"EA",x"18",x"69",x"01",x"29",x"07",x"85", -- 0x0948
    x"EA",x"85",x"EB",x"8D",x"04",x"01",x"18",x"69", -- 0x0950
    x"34",x"A2",x"34",x"A0",x"48",x"20",x"C2",x"AE", -- 0x0958
    x"20",x"59",x"AB",x"20",x"FC",x"A9",x"A6",x"A2", -- 0x0960
    x"85",x"A2",x"E0",x"01",x"F0",x"1A",x"C9",x"00", -- 0x0968
    x"F0",x"16",x"A5",x"E7",x"49",x"01",x"85",x"E7", -- 0x0970
    x"8D",x"05",x"01",x"18",x"69",x"34",x"A2",x"1C", -- 0x0978
    x"A0",x"38",x"20",x"C2",x"AE",x"20",x"59",x"AB", -- 0x0980
    x"20",x"E5",x"A9",x"F0",x"A2",x"20",x"08",x"AA", -- 0x0988
    x"AD",x"04",x"01",x"85",x"EA",x"85",x"EB",x"A9", -- 0x0990
    x"02",x"85",x"E8",x"85",x"E9",x"AE",x"05",x"01", -- 0x0998
    x"BD",x"8D",x"AB",x"85",x"E9",x"A9",x"00",x"85", -- 0x09A0
    x"E7",x"20",x"59",x"AB",x"20",x"A1",x"AE",x"A2", -- 0x09A8
    x"FF",x"9A",x"4C",x"E3",x"A0",x"A0",x"05",x"A9", -- 0x09B0
    x"F0",x"20",x"95",x"AE",x"88",x"B9",x"C6",x"A9", -- 0x09B8
    x"8D",x"0C",x"90",x"D0",x"F2",x"60",x"00",x"E3", -- 0x09C0
    x"DB",x"D6",x"D2",x"C9",x"A2",x"06",x"86",x"21", -- 0x09C8
    x"BD",x"9B",x"AB",x"48",x"BC",x"95",x"AB",x"BD", -- 0x09D0
    x"8F",x"AB",x"AA",x"68",x"20",x"4F",x"AE",x"A6", -- 0x09D8
    x"21",x"CA",x"10",x"EA",x"60",x"A9",x"EF",x"20", -- 0x09E0
    x"EB",x"AC",x"29",x"80",x"D0",x"17",x"F0",x"09", -- 0x09E8
    x"A9",x"BF",x"20",x"EB",x"AC",x"29",x"80",x"D0", -- 0x09F0
    x"0C",x"A9",x"01",x"60",x"A9",x"DF",x"20",x"EB", -- 0x09F8
    x"AC",x"29",x"80",x"F0",x"F4",x"A9",x"00",x"60", -- 0x0A00
    x"20",x"93",x"AE",x"20",x"E5",x"A9",x"D0",x"F8", -- 0x0A08
    x"60",x"20",x"A1",x"AE",x"A9",x"2F",x"8D",x"0E", -- 0x0A10
    x"90",x"A6",x"E7",x"D6",x"E8",x"30",x"25",x"20", -- 0x0A18
    x"33",x"AB",x"20",x"D1",x"AB",x"A2",x"0A",x"20", -- 0x0A20
    x"93",x"AE",x"20",x"93",x"AE",x"8A",x"48",x"29", -- 0x0A28
    x"01",x"F0",x"06",x"20",x"B2",x"AB",x"4C",x"3C", -- 0x0A30
    x"AA",x"20",x"A1",x"AB",x"68",x"AA",x"CA",x"10", -- 0x0A38
    x"E6",x"4C",x"20",x"A1",x"20",x"D1",x"AB",x"A6", -- 0x0A40
    x"E7",x"A9",x"FF",x"95",x"E8",x"A0",x"08",x"84", -- 0x0A48
    x"0E",x"A2",x"18",x"86",x"0D",x"20",x"CD",x"AD", -- 0x0A50
    x"32",x"31",x"30",x"2E",x"16",x"16",x"2D",x"2C", -- 0x0A58
    x"2E",x"2A",x"00",x"20",x"A1",x"AE",x"A9",x"32", -- 0x0A60
    x"85",x"00",x"20",x"33",x"AB",x"A2",x"0A",x"20", -- 0x0A68
    x"93",x"AE",x"CA",x"D0",x"FA",x"A2",x"18",x"86", -- 0x0A70
    x"0D",x"A0",x"08",x"84",x"0E",x"20",x"CD",x"AD", -- 0x0A78
    x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16", -- 0x0A80
    x"16",x"16",x"00",x"4C",x"22",x"AA",x"A0",x"02", -- 0x0A88
    x"A9",x"00",x"19",x"EE",x"00",x"19",x"F0",x"00", -- 0x0A90
    x"19",x"F4",x"00",x"88",x"10",x"F4",x"24",x"E8", -- 0x0A98
    x"D0",x"03",x"20",x"66",x"B0",x"A0",x"01",x"84", -- 0x0AA0
    x"0C",x"E6",x"0C",x"A5",x"0C",x"C9",x"14",x"F0", -- 0x0AA8
    x"23",x"0A",x"0A",x"0A",x"A8",x"A2",x"00",x"20", -- 0x0AB0
    x"CD",x"AD",x"16",x"16",x"16",x"16",x"16",x"16", -- 0x0AB8
    x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16", -- 0x0AC0
    x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16", -- 0x0AC8
    x"00",x"4C",x"A9",x"AA",x"A2",x"02",x"A0",x"04", -- 0x0AD0
    x"A9",x"07",x"20",x"4F",x"AE",x"20",x"59",x"AB", -- 0x0AD8
    x"A2",x"10",x"A0",x"28",x"20",x"CD",x"AD",x"1B", -- 0x0AE0
    x"34",x"26",x"24",x"22",x"31",x"2A",x"22",x"16", -- 0x0AE8
    x"32",x"31",x"30",x"2E",x"00",x"A2",x"10",x"A0", -- 0x0AF0
    x"40",x"20",x"CD",x"AD",x"1B",x"38",x"26",x"2D", -- 0x0AF8
    x"28",x"22",x"20",x"2D",x"29",x"24",x"00",x"20", -- 0x0B00
    x"70",x"AB",x"20",x"22",x"AE",x"A5",x"0C",x"F0", -- 0x0B08
    x"10",x"20",x"E5",x"A9",x"D0",x"0B",x"20",x"F0", -- 0x0B10
    x"A9",x"F0",x"EC",x"20",x"59",x"AB",x"4C",x"71", -- 0x0B18
    x"A8",x"20",x"59",x"AB",x"20",x"90",x"A9",x"A2", -- 0x0B20
    x"FF",x"9A",x"4C",x"E3",x"A0",x"A2",x"FF",x"9A", -- 0x0B28
    x"4C",x"44",x"A0",x"A5",x"E7",x"49",x"01",x"AA", -- 0x0B30
    x"B5",x"E8",x"30",x"14",x"86",x"E7",x"A2",x"1D", -- 0x0B38
    x"B5",x"C9",x"A8",x"BD",x"E1",x"1F",x"95",x"C9", -- 0x0B40
    x"98",x"9D",x"E1",x"1F",x"CA",x"10",x"F1",x"60", -- 0x0B48
    x"A6",x"E7",x"B5",x"E8",x"10",x"36",x"4C",x"8E", -- 0x0B50
    x"AA",x"A9",x"0E",x"8D",x"0F",x"90",x"A9",x"2F", -- 0x0B58
    x"8D",x"0E",x"90",x"A9",x"00",x"85",x"A9",x"85", -- 0x0B60
    x"9E",x"85",x"9F",x"A9",x"24",x"85",x"A0",x"60", -- 0x0B68
    x"E6",x"9E",x"D0",x"18",x"E6",x"9F",x"D0",x"14", -- 0x0B70
    x"A5",x"A9",x"D0",x"04",x"C6",x"A0",x"D0",x"0C", -- 0x0B78
    x"A2",x"07",x"86",x"A9",x"20",x"FF",x"AD",x"09", -- 0x0B80
    x"08",x"8D",x"0F",x"90",x"60",x"FF",x"02",x"00", -- 0x0B88
    x"01",x"02",x"07",x"08",x"0A",x"00",x"01",x"06", -- 0x0B90
    x"07",x"09",x"0A",x"07",x"06",x"07",x"0F",x"03", -- 0x0B98
    x"07",x"A2",x"38",x"A0",x"A8",x"20",x"CD",x"AD", -- 0x0BA0
    x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16", -- 0x0BA8
    x"00",x"60",x"A2",x"38",x"A0",x"A8",x"20",x"CD", -- 0x0BB0
    x"AD",x"28",x"27",x"31",x"19",x"2E",x"2A",x"00", -- 0x0BB8
    x"A2",x"54",x"A0",x"A8",x"A5",x"E7",x"18",x"69", -- 0x0BC0
    x"34",x"20",x"C2",x"AE",x"60",x"A6",x"E7",x"F6", -- 0x0BC8
    x"E8",x"20",x"B2",x"AB",x"A2",x"00",x"A0",x"A8", -- 0x0BD0
    x"20",x"CD",x"AD",x"16",x"16",x"16",x"16",x"16", -- 0x0BD8
    x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16", -- 0x0BE0
    x"16",x"00",x"A0",x"A8",x"84",x"0E",x"A2",x"00", -- 0x0BE8
    x"86",x"0D",x"A4",x"E7",x"B6",x"E8",x"86",x"A3", -- 0x0BF0
    x"30",x"2E",x"F0",x"16",x"C6",x"A3",x"E0",x"0D", -- 0x0BF8
    x"90",x"04",x"A2",x"0C",x"86",x"A3",x"A9",x"15", -- 0x0C00
    x"20",x"C6",x"AE",x"A5",x"0D",x"18",x"69",x"04", -- 0x0C08
    x"85",x"0D",x"A9",x"16",x"20",x"C6",x"AE",x"C6", -- 0x0C10
    x"A3",x"10",x"EB",x"A6",x"E7",x"B5",x"E8",x"C9", -- 0x0C18
    x"0D",x"90",x"05",x"A9",x"25",x"4C",x"C6",x"AE", -- 0x0C20
    x"60",x"20",x"A1",x"AE",x"A6",x"E7",x"A5",x"6C", -- 0x0C28
    x"C9",x"08",x"F0",x"02",x"F6",x"6C",x"F8",x"B5", -- 0x0C30
    x"EA",x"18",x"69",x"01",x"95",x"EA",x"D8",x"20", -- 0x0C38
    x"48",x"AC",x"A2",x"FF",x"9A",x"4C",x"F8",x"A0", -- 0x0C40
    x"A9",x"A0",x"85",x"0E",x"A9",x"58",x"85",x"0D", -- 0x0C48
    x"A9",x"16",x"20",x"C6",x"AE",x"A5",x"0D",x"38", -- 0x0C50
    x"E9",x"04",x"10",x"F2",x"A2",x"54",x"86",x"0D", -- 0x0C58
    x"A6",x"E7",x"B5",x"EA",x"F8",x"18",x"69",x"01", -- 0x0C60
    x"D8",x"4A",x"4A",x"4A",x"4A",x"F0",x"12",x"85", -- 0x0C68
    x"21",x"A9",x"17",x"20",x"C6",x"AE",x"A5",x"0D", -- 0x0C70
    x"38",x"E9",x"04",x"85",x"0D",x"C6",x"21",x"D0", -- 0x0C78
    x"F0",x"A6",x"E7",x"B5",x"EA",x"F8",x"18",x"69", -- 0x0C80
    x"01",x"D8",x"29",x"0F",x"F0",x"12",x"85",x"21", -- 0x0C88
    x"A9",x"18",x"20",x"C6",x"AE",x"A5",x"0D",x"38", -- 0x0C90
    x"E9",x"04",x"85",x"0D",x"C6",x"21",x"D0",x"F0", -- 0x0C98
    x"60",x"20",x"F0",x"A9",x"F0",x"03",x"4C",x"71", -- 0x0CA0
    x"A8",x"20",x"E5",x"A9",x"F0",x"09",x"20",x"90", -- 0x0CA8
    x"A9",x"A2",x"FF",x"9A",x"4C",x"E3",x"A0",x"20", -- 0x0CB0
    x"DE",x"AC",x"90",x"3A",x"A9",x"20",x"8D",x"0E", -- 0x0CB8
    x"90",x"20",x"93",x"AE",x"20",x"D8",x"AC",x"20", -- 0x0CC0
    x"70",x"AB",x"20",x"DE",x"AC",x"90",x"F8",x"20", -- 0x0CC8
    x"D8",x"AC",x"20",x"93",x"AE",x"4C",x"59",x"AB", -- 0x0CD0
    x"20",x"DE",x"AC",x"B0",x"FB",x"60",x"A9",x"EF", -- 0x0CD8
    x"20",x"EB",x"AC",x"29",x"01",x"D0",x"02",x"38", -- 0x0CE0
    x"60",x"18",x"60",x"8D",x"20",x"91",x"AD",x"21", -- 0x0CE8
    x"91",x"CD",x"21",x"91",x"D0",x"F8",x"60",x"48", -- 0x0CF0
    x"86",x"00",x"A5",x"E7",x"0A",x"18",x"65",x"E7", -- 0x0CF8
    x"AA",x"68",x"F8",x"18",x"75",x"EE",x"95",x"EE", -- 0x0D00
    x"A5",x"00",x"75",x"EF",x"95",x"EF",x"A9",x"00", -- 0x0D08
    x"75",x"F0",x"95",x"F0",x"D8",x"86",x"0C",x"A4", -- 0x0D10
    x"E7",x"B5",x"EF",x"C9",x"70",x"90",x"0E",x"B9", -- 0x0D18
    x"EC",x"00",x"D0",x"07",x"A6",x"E7",x"F6",x"EC", -- 0x0D20
    x"20",x"CD",x"AB",x"A6",x"0C",x"E8",x"E8",x"86", -- 0x0D28
    x"00",x"A0",x"02",x"B5",x"EE",x"D9",x"F4",x"00", -- 0x0D30
    x"90",x"15",x"F0",x"02",x"B0",x"04",x"CA",x"88", -- 0x0D38
    x"10",x"F1",x"A6",x"00",x"A0",x"02",x"B5",x"EE", -- 0x0D40
    x"99",x"F4",x"00",x"CA",x"88",x"10",x"F7",x"A2", -- 0x0D48
    x"20",x"A0",x"00",x"A9",x"F4",x"85",x"22",x"A9", -- 0x0D50
    x"00",x"85",x"23",x"A9",x"02",x"20",x"80",x"AD", -- 0x0D58
    x"A9",x"EE",x"85",x"22",x"A9",x"00",x"85",x"23", -- 0x0D60
    x"A2",x"00",x"A0",x"00",x"A9",x"02",x"20",x"80", -- 0x0D68
    x"AD",x"AD",x"05",x"01",x"F0",x"56",x"A9",x"F1", -- 0x0D70
    x"85",x"22",x"A2",x"40",x"A0",x"00",x"A9",x"02", -- 0x0D78
    x"86",x"0D",x"84",x"0E",x"85",x"24",x"A2",x"00", -- 0x0D80
    x"86",x"AA",x"A4",x"24",x"B1",x"22",x"48",x"4A", -- 0x0D88
    x"4A",x"4A",x"4A",x"18",x"69",x"33",x"C9",x"33", -- 0x0D90
    x"D0",x"04",x"A6",x"AA",x"F0",x"07",x"A2",x"01", -- 0x0D98
    x"86",x"AA",x"20",x"C6",x"AE",x"A5",x"0D",x"18", -- 0x0DA0
    x"69",x"04",x"85",x"0D",x"68",x"29",x"0F",x"18", -- 0x0DA8
    x"69",x"33",x"C9",x"33",x"D0",x"04",x"A6",x"AA", -- 0x0DB0
    x"F0",x"07",x"A2",x"01",x"86",x"AA",x"20",x"C6", -- 0x0DB8
    x"AE",x"A5",x"0D",x"18",x"69",x"04",x"85",x"0D", -- 0x0DC0
    x"C6",x"24",x"10",x"BE",x"60",x"86",x"0D",x"84", -- 0x0DC8
    x"0E",x"68",x"85",x"2C",x"68",x"85",x"2D",x"D0", -- 0x0DD0
    x"10",x"A0",x"00",x"B1",x"2C",x"F0",x"12",x"20", -- 0x0DD8
    x"C6",x"AE",x"A5",x"0D",x"18",x"69",x"04",x"85", -- 0x0DE0
    x"0D",x"E6",x"2C",x"D0",x"EC",x"E6",x"2D",x"D0", -- 0x0DE8
    x"E8",x"A5",x"2D",x"48",x"A5",x"2C",x"48",x"60", -- 0x0DF0
    x"A5",x"0C",x"29",x"10",x"D0",x"FA",x"60",x"AD", -- 0x0DF8
    x"04",x"90",x"6D",x"01",x"01",x"EE",x"03",x"01", -- 0x0E00
    x"EE",x"00",x"01",x"AC",x"03",x"01",x"71",x"FF", -- 0x0E08
    x"6D",x"04",x"90",x"8D",x"01",x"01",x"3D",x"1A", -- 0x0E10
    x"AE",x"60",x"01",x"03",x"07",x"0F",x"1F",x"3F", -- 0x0E18
    x"7F",x"FF",x"A0",x"03",x"A9",x"FF",x"C0",x"02", -- 0x0E20
    x"F0",x"09",x"8D",x"22",x"91",x"AD",x"11",x"91", -- 0x0E28
    x"4C",x"3A",x"AE",x"4A",x"8D",x"22",x"91",x"AD", -- 0x0E30
    x"20",x"91",x"39",x"4B",x"AE",x"99",x"08",x"00", -- 0x0E38
    x"88",x"10",x"E1",x"AD",x"11",x"91",x"29",x"20", -- 0x0E40
    x"85",x"0C",x"60",x"10",x"04",x"80",x"08",x"86", -- 0x0E48
    x"06",x"84",x"07",x"48",x"20",x"8A",x"AE",x"A0", -- 0x0E50
    x"15",x"68",x"91",x"04",x"88",x"10",x"FB",x"A4", -- 0x0E58
    x"07",x"C4",x"06",x"F0",x"24",x"88",x"10",x"E9", -- 0x0E60
    x"A9",x"10",x"85",x"03",x"A9",x"00",x"85",x"02", -- 0x0E68
    x"A8",x"A2",x"0F",x"91",x"02",x"99",x"20",x"1E", -- 0x0E70
    x"C8",x"D0",x"F8",x"E6",x"03",x"CA",x"D0",x"F3", -- 0x0E78
    x"60",x"B1",x"F7",x"85",x"02",x"B1",x"F9",x"85", -- 0x0E80
    x"03",x"60",x"B1",x"FB",x"85",x"04",x"B1",x"FD", -- 0x0E88
    x"85",x"05",x"60",x"A9",x"FF",x"38",x"48",x"E9", -- 0x0E90
    x"01",x"D0",x"FC",x"68",x"E9",x"01",x"D0",x"F6", -- 0x0E98
    x"60",x"20",x"B0",x"AE",x"20",x"B6",x"AE",x"20", -- 0x0EA0
    x"BC",x"AE",x"A9",x"00",x"8D",x"0D",x"90",x"60", -- 0x0EA8
    x"A9",x"00",x"8D",x"0A",x"90",x"60",x"A9",x"00", -- 0x0EB0
    x"8D",x"0B",x"90",x"60",x"A9",x"00",x"8D",x"0C", -- 0x0EB8
    x"90",x"60",x"86",x"0D",x"84",x"0E",x"A6",x"0D", -- 0x0EC0
    x"85",x"18",x"8A",x"29",x"03",x"85",x"19",x"8A", -- 0x0EC8
    x"4A",x"4A",x"85",x"14",x"A5",x"18",x"0A",x"A8", -- 0x0ED0
    x"B9",x"E4",x"B1",x"85",x"1A",x"C8",x"B9",x"E4", -- 0x0ED8
    x"B1",x"85",x"1B",x"A0",x"00",x"B1",x"1A",x"85", -- 0x0EE0
    x"11",x"C8",x"B1",x"1A",x"85",x"12",x"A5",x"1A", -- 0x0EE8
    x"18",x"69",x"02",x"85",x"15",x"A5",x"1B",x"69", -- 0x0EF0
    x"00",x"85",x"16",x"A9",x"00",x"85",x"1C",x"A5", -- 0x0EF8
    x"12",x"85",x"17",x"A5",x"0E",x"85",x"1D",x"A4", -- 0x0F00
    x"14",x"C0",x"16",x"B0",x"4A",x"20",x"81",x"AE", -- 0x0F08
    x"A5",x"17",x"C5",x"12",x"F0",x"42",x"C9",x"01", -- 0x0F10
    x"F0",x"42",x"A2",x"04",x"A4",x"11",x"84",x"13", -- 0x0F18
    x"A9",x"00",x"A4",x"1C",x"20",x"6D",x"AF",x"A4", -- 0x0F20
    x"1D",x"48",x"AD",x"02",x"01",x"F0",x"08",x"10", -- 0x0F28
    x"0C",x"68",x"31",x"02",x"4C",x"47",x"AF",x"68", -- 0x0F30
    x"11",x"02",x"4C",x"47",x"AF",x"B1",x"02",x"3D", -- 0x0F38
    x"64",x"AF",x"85",x"00",x"68",x"05",x"00",x"91", -- 0x0F40
    x"02",x"E6",x"1C",x"E6",x"1D",x"C6",x"13",x"D0", -- 0x0F48
    x"CF",x"E6",x"14",x"C6",x"17",x"D0",x"AC",x"60", -- 0x0F50
    x"A6",x"19",x"10",x"C0",x"A9",x"05",x"18",x"65", -- 0x0F58
    x"19",x"AA",x"D0",x"B8",x"00",x"C0",x"F0",x"FC", -- 0x0F60
    x"00",x"FF",x"3F",x"0F",x"03",x"85",x"0F",x"86", -- 0x0F68
    x"10",x"E0",x"04",x"90",x"1B",x"F0",x"21",x"98", -- 0x0F70
    x"38",x"E5",x"11",x"A8",x"B1",x"15",x"A8",x"A5", -- 0x0F78
    x"19",x"18",x"69",x"FC",x"AA",x"98",x"0A",x"0A", -- 0x0F80
    x"E8",x"D0",x"FB",x"05",x"0F",x"A6",x"10",x"60", -- 0x0F88
    x"B1",x"15",x"20",x"A4",x"AF",x"4C",x"8B",x"AF", -- 0x0F90
    x"B1",x"15",x"20",x"A4",x"AF",x"05",x"0F",x"85", -- 0x0F98
    x"0F",x"4C",x"77",x"AF",x"A6",x"19",x"F0",x"05", -- 0x0FA0
    x"4A",x"4A",x"CA",x"D0",x"FB",x"60",x"00",x"0A", -- 0x0FA8
    x"0C",x"0F",x"0E",x"0D",x"0E",x"0D",x"0C",x"0D", -- 0x0FB0
    x"0C",x"0B",x"00",x"00",x"00",x"01",x"01",x"02", -- 0x0FB8
    x"02",x"07",x"00",x"00",x"90",x"40",x"40",x"40", -- 0x0FC0
    x"40",x"40",x"00",x"1A",x"19",x"1B",x"00",x"17", -- 0x0FC8
    x"18",x"16",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FD8
    x"00",x"00",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x0FE0
    x"04",x"04",x"04",x"04",x"04",x"04",x"06",x"06", -- 0x0FE8
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0FF0
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0FF8
    x"40",x"40",x"40",x"40",x"40",x"40",x"50",x"50", -- 0x1000
    x"50",x"50",x"50",x"50",x"60",x"60",x"2D",x"27", -- 0x1008
    x"21",x"1B",x"15",x"0F",x"09",x"03",x"2D",x"27", -- 0x1010
    x"21",x"1B",x"15",x"0F",x"09",x"03",x"27",x"21", -- 0x1018
    x"1B",x"15",x"0F",x"09",x"27",x"21",x"1B",x"15", -- 0x1020
    x"0F",x"09",x"0F",x"21",x"3C",x"3C",x"3C",x"3C", -- 0x1028
    x"3C",x"3C",x"3C",x"3C",x"32",x"32",x"32",x"32", -- 0x1030
    x"32",x"32",x"32",x"32",x"28",x"28",x"28",x"28", -- 0x1038
    x"28",x"28",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E", -- 0x1040
    x"14",x"14",x"19",x"18",x"13",x"12",x"0C",x"0B", -- 0x1048
    x"04",x"03",x"1A",x"17",x"14",x"11",x"0D",x"0A", -- 0x1050
    x"05",x"02",x"1B",x"16",x"15",x"10",x"0E",x"09", -- 0x1058
    x"06",x"01",x"0F",x"08",x"07",x"00",x"A2",x"1C", -- 0x1060
    x"A0",x"00",x"20",x"CD",x"AD",x"22",x"1E",x"2E", -- 0x1068
    x"16",x"2F",x"2E",x"2A",x"2B",x"00",x"60",x"07", -- 0x1070
    x"06",x"05",x"04",x"03",x"02",x"02",x"01",x"01", -- 0x1078
    x"05",x"05",x"06",x"06",x"07",x"08",x"09",x"0A", -- 0x1080
    x"0B",x"11",x"20",x"20",x"2C",x"10",x"C0",x"B0", -- 0x1088
    x"D2",x"B0",x"F3",x"B0",x"14",x"B1",x"41",x"B1", -- 0x1090
    x"52",x"B1",x"64",x"B1",x"85",x"B1",x"A6",x"B1", -- 0x1098
    x"D3",x"B1",x"80",x"80",x"80",x"80",x"00",x"00", -- 0x10A0
    x"00",x"00",x"80",x"80",x"80",x"80",x"00",x"00", -- 0x10A8
    x"00",x"00",x"80",x"80",x"80",x"00",x"00",x"00", -- 0x10B0
    x"80",x"80",x"80",x"00",x"00",x"00",x"00",x"80", -- 0x10B8
    x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00", -- 0x10C0
    x"00",x"01",x"00",x"01",x"01",x"01",x"01",x"01", -- 0x10C8
    x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00", -- 0x10D0
    x"00",x"00",x"01",x"00",x"00",x"01",x"00",x"00", -- 0x10D8
    x"00",x"01",x"00",x"00",x"01",x"01",x"00",x"01", -- 0x10E0
    x"00",x"01",x"01",x"00",x"01",x"01",x"01",x"01", -- 0x10E8
    x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"00", -- 0x10F0
    x"01",x"00",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x10F8
    x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x1100
    x"00",x"01",x"01",x"01",x"00",x"01",x"01",x"01", -- 0x1108
    x"00",x"01",x"01",x"00",x"00",x"01",x"00",x"01", -- 0x1110
    x"01",x"00",x"01",x"01",x"00",x"01",x"01",x"01", -- 0x1118
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x1120
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x1128
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x1130
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x1138
    x"00",x"00",x"00",x"00",x"01",x"00",x"01",x"01", -- 0x1140
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00", -- 0x1148
    x"01",x"00",x"00",x"01",x"01",x"01",x"01",x"01", -- 0x1150
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF", -- 0x1158
    x"FF",x"FF",x"FF",x"FF",x"00",x"02",x"02",x"02", -- 0x1160
    x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x1168
    x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x1170
    x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x1178
    x"02",x"02",x"02",x"02",x"02",x"00",x"02",x"02", -- 0x1180
    x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x1188
    x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x1190
    x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x1198
    x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"02", -- 0x11A0
    x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x11A8
    x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01", -- 0x11B0
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x11B8
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x11C0
    x"01",x"01",x"02",x"01",x"01",x"02",x"02",x"02", -- 0x11C8
    x"02",x"02",x"02",x"00",x"02",x"02",x"02",x"02", -- 0x11D0
    x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x11D8
    x"02",x"02",x"02",x"02",x"5E",x"B2",x"72",x"B2", -- 0x11E0
    x"86",x"B2",x"9C",x"B2",x"B2",x"B2",x"C6",x"B2", -- 0x11E8
    x"DA",x"B2",x"EE",x"B2",x"02",x"B3",x"16",x"B3", -- 0x11F0
    x"2A",x"B3",x"40",x"B3",x"52",x"B3",x"64",x"B3", -- 0x11F8
    x"76",x"B3",x"88",x"B3",x"9A",x"B3",x"AC",x"B3", -- 0x1200
    x"BE",x"B3",x"C4",x"B3",x"C9",x"B3",x"CD",x"B3", -- 0x1208
    x"D7",x"B3",x"E1",x"B3",x"EB",x"B3",x"F5",x"B3", -- 0x1210
    x"FF",x"B3",x"09",x"B4",x"13",x"B4",x"1D",x"B4", -- 0x1218
    x"27",x"B4",x"31",x"B4",x"3B",x"B4",x"45",x"B4", -- 0x1220
    x"4F",x"B4",x"59",x"B4",x"63",x"B4",x"6D",x"B4", -- 0x1228
    x"77",x"B4",x"81",x"B4",x"8B",x"B4",x"95",x"B4", -- 0x1230
    x"9F",x"B4",x"A9",x"B4",x"B3",x"B4",x"BD",x"B4", -- 0x1238
    x"C7",x"B4",x"D1",x"B4",x"DB",x"B4",x"E5",x"B4", -- 0x1240
    x"EF",x"B4",x"F9",x"B4",x"03",x"B5",x"0D",x"B5", -- 0x1248
    x"17",x"B5",x"21",x"B5",x"2B",x"B5",x"35",x"B5", -- 0x1250
    x"3F",x"B5",x"49",x"B5",x"53",x"B5",x"09",x"03", -- 0x1258
    x"00",x"00",x"04",x"01",x"0D",x"01",x"05",x"0C", -- 0x1260
    x"00",x"00",x"00",x"10",x"40",x"70",x"40",x"50", -- 0x1268
    x"30",x"00",x"09",x"03",x"00",x"00",x"00",x"04", -- 0x1270
    x"01",x"0D",x"01",x"0C",x"00",x"00",x"00",x"00", -- 0x1278
    x"10",x"40",x"70",x"40",x"30",x"00",x"0A",x"03", -- 0x1280
    x"00",x"00",x"00",x"08",x"01",x"0D",x"01",x"0B", -- 0x1288
    x"0C",x"00",x"00",x"00",x"00",x"20",x"40",x"70", -- 0x1290
    x"40",x"E0",x"30",x"00",x"0A",x"03",x"00",x"00", -- 0x1298
    x"00",x"00",x"08",x"01",x"0D",x"03",x"08",x"00", -- 0x12A0
    x"00",x"00",x"00",x"00",x"20",x"40",x"70",x"C0", -- 0x12A8
    x"20",x"00",x"09",x"03",x"00",x"00",x"09",x"0E", -- 0x12B0
    x"0F",x"03",x"03",x"00",x"00",x"00",x"00",x"10", -- 0x12B8
    x"60",x"B0",x"C0",x"C0",x"C0",x"00",x"09",x"03", -- 0x12C0
    x"00",x"00",x"00",x"04",x"08",x"0E",x"03",x"03", -- 0x12C8
    x"00",x"00",x"00",x"00",x"10",x"B0",x"F0",x"C0", -- 0x12D0
    x"C0",x"00",x"09",x"03",x"00",x"00",x"0D",x"0B", -- 0x12D8
    x"0A",x"02",x"02",x"00",x"00",x"00",x"00",x"10", -- 0x12E0
    x"70",x"E0",x"80",x"80",x"80",x"00",x"09",x"03", -- 0x12E8
    x"00",x"00",x"00",x"04",x"0C",x"0B",x"02",x"02", -- 0x12F0
    x"00",x"00",x"00",x"00",x"10",x"E0",x"A0",x"80", -- 0x12F8
    x"80",x"00",x"09",x"03",x"00",x"00",x"02",x"09", -- 0x1300
    x"11",x"20",x"01",x"18",x"00",x"00",x"00",x"B0", -- 0x1308
    x"14",x"40",x"C8",x"20",x"C0",x"00",x"09",x"03", -- 0x1310
    x"00",x"00",x"02",x"21",x"18",x"22",x"28",x"13", -- 0x1318
    x"08",x"00",x"60",x"A0",x"18",x"48",x"88",x"10", -- 0x1320
    x"20",x"40",x"0A",x"03",x"00",x"00",x"00",x"00", -- 0x1328
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1330
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1338
    x"08",x"03",x"00",x"28",x"2F",x"0D",x"0D",x"2F", -- 0x1340
    x"28",x"00",x"00",x"A0",x"E0",x"C0",x"C0",x"E0", -- 0x1348
    x"A0",x"00",x"08",x"03",x"00",x"23",x"0B",x"3D", -- 0x1350
    x"3D",x"0B",x"23",x"00",x"00",x"20",x"80",x"F0", -- 0x1358
    x"F0",x"80",x"20",x"00",x"08",x"03",x"00",x"02", -- 0x1360
    x"38",x"0D",x"29",x"0C",x"2E",x"00",x"00",x"E0", -- 0x1368
    x"C0",x"A0",x"C0",x"B0",x"00",x"00",x"08",x"03", -- 0x1370
    x"3C",x"8E",x"AC",x"A9",x"2D",x"EF",x"C3",x"0F", -- 0x1378
    x"A0",x"B0",x"B8",x"F8",x"B8",x"B0",x"80",x"A0", -- 0x1380
    x"08",x"03",x"0F",x"2B",x"E3",x"E1",x"E1",x"E3", -- 0x1388
    x"2B",x"0F",x"C0",x"A0",x"2C",x"2C",x"2C",x"2C", -- 0x1390
    x"A0",x"C0",x"08",x"03",x"02",x"02",x"0F",x"0F", -- 0x1398
    x"12",x"1E",x"1E",x"12",x"00",x"00",x"C0",x"C0", -- 0x13A0
    x"10",x"D0",x"D0",x"10",x"08",x"03",x"00",x"00", -- 0x13A8
    x"0F",x"0F",x"12",x"1E",x"1E",x"12",x"00",x"00", -- 0x13B0
    x"C0",x"C0",x"10",x"D0",x"D0",x"10",x"04",x"01", -- 0x13B8
    x"80",x"80",x"80",x"00",x"03",x"01",x"00",x"00", -- 0x13C0
    x"00",x"02",x"01",x"C0",x"C0",x"08",x"01",x"00", -- 0x13C8
    x"00",x"18",x"5A",x"66",x"5A",x"66",x"00",x"08", -- 0x13D0
    x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13D8
    x"00",x"08",x"01",x"00",x"7E",x"7E",x"7E",x"7E", -- 0x13E0
    x"60",x"60",x"60",x"08",x"01",x"00",x"00",x"7C", -- 0x13E8
    x"7C",x"7C",x"40",x"40",x"40",x"08",x"01",x"66", -- 0x13F0
    x"66",x"66",x"3C",x"18",x"18",x"18",x"00",x"08", -- 0x13F8
    x"01",x"7C",x"66",x"66",x"7C",x"66",x"66",x"7C", -- 0x1400
    x"00",x"08",x"01",x"3C",x"66",x"60",x"7C",x"60", -- 0x1408
    x"60",x"60",x"00",x"08",x"01",x"66",x"66",x"3C", -- 0x1410
    x"18",x"3C",x"66",x"66",x"00",x"08",x"01",x"66", -- 0x1418
    x"66",x"66",x"66",x"66",x"66",x"3C",x"00",x"08", -- 0x1420
    x"01",x"66",x"66",x"66",x"7E",x"66",x"66",x"66", -- 0x1428
    x"00",x"08",x"01",x"3C",x"66",x"60",x"60",x"60", -- 0x1430
    x"66",x"3C",x"00",x"08",x"01",x"7E",x"18",x"18", -- 0x1438
    x"18",x"18",x"18",x"7E",x"00",x"08",x"01",x"7C", -- 0x1440
    x"66",x"66",x"66",x"66",x"66",x"7C",x"00",x"08", -- 0x1448
    x"01",x"7E",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x1450
    x"00",x"08",x"01",x"3C",x"42",x"9D",x"A1",x"A1", -- 0x1458
    x"9D",x"42",x"3C",x"08",x"01",x"3C",x"66",x"60", -- 0x1460
    x"3C",x"06",x"66",x"3C",x"00",x"08",x"01",x"00", -- 0x1468
    x"00",x"10",x"10",x"7C",x"10",x"10",x"00",x"08", -- 0x1470
    x"01",x"00",x"00",x"00",x"7E",x"7E",x"00",x"00", -- 0x1478
    x"00",x"08",x"01",x"60",x"60",x"60",x"60",x"60", -- 0x1480
    x"60",x"7E",x"00",x"08",x"01",x"7C",x"66",x"66", -- 0x1488
    x"7C",x"60",x"60",x"60",x"00",x"08",x"01",x"66", -- 0x1490
    x"66",x"76",x"6E",x"66",x"66",x"66",x"00",x"08", -- 0x1498
    x"01",x"7C",x"66",x"66",x"7C",x"78",x"6C",x"66", -- 0x14A0
    x"00",x"08",x"01",x"66",x"6C",x"78",x"70",x"78", -- 0x14A8
    x"6C",x"66",x"00",x"08",x"01",x"66",x"66",x"66", -- 0x14B0
    x"66",x"66",x"3C",x"18",x"00",x"08",x"01",x"3C", -- 0x14B8
    x"66",x"66",x"66",x"66",x"66",x"3C",x"00",x"08", -- 0x14C0
    x"01",x"3C",x"66",x"60",x"7C",x"60",x"66",x"3C", -- 0x14C8
    x"00",x"08",x"01",x"3E",x"0C",x"0C",x"0C",x"0C", -- 0x14D0
    x"6C",x"38",x"00",x"08",x"01",x"66",x"7E",x"66", -- 0x14D8
    x"66",x"66",x"66",x"66",x"00",x"08",x"01",x"3C", -- 0x14E0
    x"66",x"66",x"7E",x"66",x"66",x"66",x"00",x"08", -- 0x14E8
    x"01",x"3C",x"66",x"60",x"6E",x"66",x"66",x"3C", -- 0x14F0
    x"00",x"08",x"01",x"3C",x"66",x"6E",x"7E",x"76", -- 0x14F8
    x"66",x"3C",x"00",x"08",x"01",x"18",x"38",x"78", -- 0x1500
    x"18",x"18",x"18",x"7E",x"00",x"08",x"01",x"3C", -- 0x1508
    x"66",x"06",x"0C",x"18",x"30",x"7E",x"00",x"08", -- 0x1510
    x"01",x"3C",x"66",x"06",x"1C",x"06",x"66",x"3C", -- 0x1518
    x"00",x"08",x"01",x"0E",x"1E",x"36",x"66",x"7E", -- 0x1520
    x"06",x"06",x"00",x"08",x"01",x"7E",x"60",x"60", -- 0x1528
    x"7C",x"06",x"66",x"3C",x"00",x"08",x"01",x"1C", -- 0x1530
    x"30",x"60",x"7C",x"66",x"66",x"3C",x"00",x"08", -- 0x1538
    x"01",x"7E",x"66",x"0C",x"18",x"18",x"18",x"18", -- 0x1540
    x"00",x"08",x"01",x"3C",x"66",x"66",x"3C",x"66", -- 0x1548
    x"66",x"3C",x"00",x"08",x"01",x"3C",x"66",x"66", -- 0x1550
    x"3E",x"06",x"0C",x"18",x"00",x"EA",x"00",x"EA", -- 0x1558
    x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x1560
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1568
    x"B0",x"99",x"6E",x"00",x"60",x"A2",x"00",x"20", -- 0x1570
    x"FF",x"AD",x"18",x"69",x"1C",x"A8",x"A2",x"08", -- 0x1578
    x"B9",x"C9",x"00",x"F0",x"B7",x"B5",x"8C",x"D0", -- 0x1580
    x"B3",x"A9",x"01",x"85",x"9A",x"86",x"95",x"84", -- 0x1588
    x"96",x"20",x"63",x"A5",x"A5",x"96",x"38",x"E9", -- 0x1590
    x"1C",x"AA",x"A0",x"07",x"84",x"95",x"0A",x"0A", -- 0x1598
    x"09",x"03",x"85",x"00",x"A9",x"02",x"85",x"01", -- 0x15A0
    x"A6",x"00",x"BC",x"CA",x"AF",x"F0",x"C5",x"B9", -- 0x15A8
    x"C9",x"00",x"F0",x"17",x"B9",x"6E",x"00",x"D0", -- 0x15B0
    x"12",x"A6",x"95",x"B5",x"8C",x"D0",x"0C",x"20", -- 0x15B8
    x"63",x"A5",x"A5",x"9A",x"0A",x"85",x"9A",x"C6", -- 0x15C0
    x"95",x"C6",x"01",x"A5",x"01",x"F0",x"A5",x"C6", -- 0x15C8
    x"00",x"10",x"D5",x"A5",x"9B",x"F0",x"9D",x"C6", -- 0x15D0
    x"9B",x"D0",x"99",x"A2",x"28",x"86",x"0D",x"A0", -- 0x15D8
    x"A8",x"84",x"0E",x"A9",x"16",x"20",x"C6",x"AE", -- 0x15E0
    x"A5",x"0D",x"38",x"E9",x"04",x"C9",x"18",x"F0", -- 0x15E8
    x"83",x"85",x"0D",x"10",x"EE",x"A5",x"9C",x"D0", -- 0x15F0
    x"57",x"C6",x"26",x"10",x"52",x"A9",x"05",x"85", -- 0x15F8
    x"26",x"20",x"22",x"AE",x"A5",x"25",x"A6",x"0A", -- 0x1600
    x"F0",x"0B",x"A6",x"08",x"D0",x"10",x"38",x"E9", -- 0x1608
    x"01",x"10",x"09",x"30",x"09",x"18",x"69",x"01", -- 0x1610
    x"C9",x"52",x"F0",x"02",x"85",x"25",x"A5",x"2B", -- 0x1618
    x"D0",x"1D",x"A5",x"0C",x"F0",x"06",x"A9",x"00", -- 0x1620
    x"85",x"6D",x"F0",x"13",x"A5",x"6D",x"D0",x"0F", -- 0x1628
    x"E6",x"6D",x"A5",x"25",x"18",x"69",x"03",x"85", -- 0x1630
    x"29",x"85",x"2B",x"A9",x"98",x"85",x"2A",x"A0", -- 0x1638
    x"98",x"A6",x"25",x"A5",x"2B",x"F0",x"03",x"A9", -- 0x1640
    x"11",x"2C",x"A9",x"10",x"4C",x"C2",x"AE",x"60", -- 0x1648
    x"C6",x"9D",x"10",x"FB",x"A9",x"0F",x"85",x"9D", -- 0x1650
    x"A2",x"07",x"20",x"FF",x"AD",x"8D",x"0D",x"90", -- 0x1658
    x"20",x"FF",x"AD",x"8D",x"0A",x"90",x"CE",x"0E", -- 0x1660
    x"90",x"A6",x"9C",x"BD",x"AE",x"AF",x"A6",x"25", -- 0x1668
    x"A0",x"98",x"20",x"C2",x"AE",x"C6",x"9C",x"D0", -- 0x1670
    x"D6",x"4C",x"11",x"AA",x"20",x"8B",x"A6",x"20", -- 0x1678
    x"8B",x"A6",x"20",x"8B",x"A6",x"20",x"8B",x"A6", -- 0x1680
    x"4C",x"BD",x"A3",x"A5",x"2B",x"F0",x"C0",x"C6", -- 0x1688
    x"28",x"10",x"BC",x"A9",x"01",x"85",x"28",x"A5", -- 0x1690
    x"2A",x"4A",x"18",x"69",x"AF",x"8D",x"0B",x"90", -- 0x1698
    x"A5",x"29",x"85",x"0D",x"A5",x"2A",x"85",x"0E", -- 0x16A0
    x"38",x"E9",x"01",x"C9",x"0F",x"F0",x"09",x"85", -- 0x16A8
    x"2A",x"85",x"0E",x"A9",x"12",x"4C",x"C6",x"AE", -- 0x16B0
    x"20",x"B6",x"AE",x"85",x"2B",x"A6",x"29",x"A4", -- 0x16B8
    x"2A",x"F0",x"8C",x"A9",x"13",x"4C",x"C2",x"AE", -- 0x16C0
    x"A6",x"E7",x"B4",x"6C",x"BE",x"77",x"B0",x"CA", -- 0x16C8
    x"20",x"FF",x"AD",x"D0",x"0E",x"A6",x"E7",x"B4", -- 0x16D0
    x"6C",x"BE",x"80",x"B0",x"B5",x"47",x"F0",x"04", -- 0x16D8
    x"CA",x"10",x"F9",x"60",x"86",x"2E",x"A4",x"96", -- 0x16E0
    x"B9",x"C9",x"00",x"F0",x"F6",x"C9",x"7C",x"B0", -- 0x16E8
    x"F2",x"18",x"69",x"0C",x"95",x"3B",x"85",x"0E", -- 0x16F0
    x"B9",x"AB",x"00",x"18",x"69",x"03",x"C9",x"54", -- 0x16F8
    x"B0",x"E1",x"95",x"2F",x"85",x"0D",x"A6",x"96", -- 0x1700
    x"A0",x"01",x"B5",x"AB",x"C5",x"25",x"90",x"07", -- 0x1708
    x"98",x"49",x"FF",x"18",x"69",x"01",x"A8",x"A6", -- 0x1710
    x"2E",x"94",x"47",x"A9",x"14",x"4C",x"C6",x"AE", -- 0x1718
    x"C6",x"A8",x"10",x"BF",x"A9",x"01",x"85",x"A8", -- 0x1720
    x"A6",x"E7",x"B4",x"6C",x"BE",x"80",x"B0",x"86", -- 0x1728
    x"2E",x"B5",x"47",x"F0",x"47",x"B5",x"3B",x"85", -- 0x1730
    x"0E",x"B5",x"2F",x"85",x"0D",x"A9",x"13",x"20", -- 0x1738
    x"C6",x"AE",x"A6",x"2E",x"B5",x"2F",x"30",x"47", -- 0x1740
    x"C9",x"54",x"B0",x"43",x"85",x"0D",x"B5",x"3B", -- 0x1748
    x"18",x"69",x"05",x"C9",x"9C",x"B0",x"38",x"95", -- 0x1750
    x"3B",x"85",x"0E",x"4A",x"85",x"00",x"A9",x"C8", -- 0x1758
    x"38",x"E5",x"00",x"8D",x"0C",x"90",x"A9",x"14", -- 0x1760
    x"20",x"C6",x"AE",x"A6",x"2E",x"B5",x"3B",x"C9", -- 0x1768
    x"93",x"90",x"09",x"B5",x"2F",x"38",x"E5",x"25", -- 0x1770
    x"C9",x"05",x"90",x"06",x"A6",x"2E",x"CA",x"10", -- 0x1778
    x"AE",x"60",x"A9",x"13",x"20",x"C6",x"AE",x"A5", -- 0x1780
    x"9C",x"D0",x"04",x"A9",x"06",x"85",x"9C",x"A6", -- 0x1788
    x"2E",x"20",x"BC",x"AE",x"95",x"47",x"F0",x"E4", -- 0x1790
    x"A9",x"10",x"4C",x"95",x"AE",x"20",x"59",x"AB", -- 0x1798
    x"20",x"68",x"AE",x"20",x"A1",x"AE",x"8D",x"02", -- 0x17A0
    x"01",x"20",x"CC",x"A9",x"A2",x"08",x"A0",x"08", -- 0x17A8
    x"20",x"CD",x"AD",x"31",x"22",x"31",x"2A",x"20", -- 0x17B0
    x"24",x"2D",x"1B",x"22",x"16",x"28",x"2A",x"2E", -- 0x17B8
    x"24",x"2E",x"29",x"22",x"24",x"00",x"A2",x"1C", -- 0x17C0
    x"A0",x"18",x"20",x"CD",x"AD",x"32",x"31",x"27", -- 0x17C8
    x"31",x"1C",x"20",x"31",x"29",x"00",x"A2",x"18", -- 0x17D0
    x"A0",x"30",x"20",x"CD",x"AD",x"28",x"2A",x"2E", -- 0x17D8
    x"24",x"24",x"16",x"1B",x"34",x"00",x"A2",x"14", -- 0x17E0
    x"A0",x"38",x"20",x"CD",x"AD",x"1B",x"2D",x"2A", -- 0x17E8
    x"16",x"2D",x"28",x"22",x"20",x"2D",x"29",x"24", -- 0x17F0
    x"00",x"A2",x"04",x"A0",x"08",x"A9",x"0F",x"20", -- 0x17F8
    x"4F",x"AE",x"A2",x"1D",x"86",x"20",x"BD",x"2C", -- 0x1800
    x"B0",x"18",x"69",x"3C",x"95",x"C9",x"BD",x"0E", -- 0x1808
    x"B0",x"95",x"AB",x"CA",x"10",x"F0",x"A9",x"15", -- 0x1810
    x"85",x"1F",x"A9",x"01",x"85",x"1E",x"20",x"85", -- 0x1818
    x"A1",x"A5",x"20",x"C9",x"1D",x"D0",x"F7",x"A2", -- 0x1820
    x"14",x"A0",x"A0",x"20",x"CD",x"AD",x"23",x"34", -- 0x1828
    x"3C",x"3B",x"36",x"16",x"31",x"22",x"31",x"2A", -- 0x1830
    x"20",x"00",x"A2",x"04",x"A0",x"A8",x"20",x"CD", -- 0x1838
    x"AD",x"31",x"27",x"27",x"16",x"2A",x"20",x"32", -- 0x1840
    x"1E",x"22",x"24",x"16",x"2A",x"2E",x"24",x"2E", -- 0x1848
    x"2A",x"2C",x"2E",x"21",x"16",x"16",x"00",x"A9", -- 0x1850
    x"01",x"8D",x"02",x"01",x"20",x"70",x"AB",x"20", -- 0x1858
    x"E5",x"A9",x"D0",x"0D",x"20",x"22",x"AE",x"A5", -- 0x1860
    x"0C",x"D0",x"F1",x"20",x"59",x"AB",x"4C",x"90", -- 0x1868
    x"A9",x"20",x"A1",x"AE",x"20",x"59",x"AB",x"20", -- 0x1870
    x"08",x"AA",x"20",x"68",x"AE",x"20",x"CC",x"A9", -- 0x1878
    x"A9",x"00",x"8D",x"02",x"01",x"20",x"4F",x"AD", -- 0x1880
    x"A2",x"10",x"A0",x"28",x"20",x"CD",x"AD",x"1B", -- 0x1888
    x"34",x"26",x"24",x"22",x"31",x"2A",x"22",x"16", -- 0x1890
    x"32",x"31",x"30",x"2E",x"00",x"A2",x"10",x"A0", -- 0x1898
    x"38",x"20",x"CD",x"AD",x"1B",x"36",x"26",x"16", -- 0x18A0
    x"16",x"28",x"27",x"31",x"19",x"2E",x"2A",x"00", -- 0x18A8
    x"AD",x"05",x"01",x"85",x"E7",x"18",x"69",x"34", -- 0x18B0
    x"A2",x"1C",x"A0",x"38",x"20",x"C2",x"AE",x"A2", -- 0x18B8
    x"10",x"A0",x"48",x"20",x"CD",x"AD",x"1B",x"38", -- 0x18C0
    x"26",x"27",x"2E",x"2C",x"2E",x"27",x"00",x"AD", -- 0x18C8
    x"04",x"01",x"85",x"EA",x"85",x"EB",x"18",x"69", -- 0x18D0
    x"34",x"A2",x"34",x"A0",x"48",x"20",x"C2",x"AE", -- 0x18D8
    x"A2",x"10",x"A0",x"70",x"20",x"CD",x"AD",x"06", -- 0x18E0
    x"16",x"16",x"16",x"16",x"16",x"04",x"16",x"16", -- 0x18E8
    x"16",x"02",x"16",x"16",x"16",x"01",x"00",x"A2", -- 0x18F0
    x"10",x"A0",x"80",x"20",x"CD",x"AD",x"39",x"33", -- 0x18F8
    x"16",x"16",x"16",x"16",x"38",x"33",x"16",x"16", -- 0x1900
    x"37",x"33",x"16",x"16",x"36",x"33",x"00",x"A2", -- 0x1908
    x"04",x"A0",x"90",x"20",x"CD",x"AD",x"34",x"38", -- 0x1910
    x"33",x"26",x"3B",x"33",x"33",x"16",x"34",x"33", -- 0x1918
    x"33",x"16",x"16",x"3B",x"33",x"16",x"16",x"39", -- 0x1920
    x"33",x"00",x"A9",x"01",x"8D",x"02",x"01",x"20", -- 0x1928
    x"70",x"AB",x"20",x"22",x"AE",x"A5",x"0C",x"F0", -- 0x1930
    x"57",x"20",x"F0",x"A9",x"A6",x"A1",x"85",x"A1", -- 0x1938
    x"E0",x"01",x"F0",x"1F",x"C9",x"00",x"F0",x"1B", -- 0x1940
    x"A5",x"EA",x"18",x"69",x"01",x"29",x"07",x"85", -- 0x1948
    x"EA",x"85",x"EB",x"8D",x"04",x"01",x"18",x"69", -- 0x1950
    x"34",x"A2",x"34",x"A0",x"48",x"20",x"C2",x"AE", -- 0x1958
    x"20",x"59",x"AB",x"20",x"FC",x"A9",x"A6",x"A2", -- 0x1960
    x"85",x"A2",x"E0",x"01",x"F0",x"1A",x"C9",x"00", -- 0x1968
    x"F0",x"16",x"A5",x"E7",x"49",x"01",x"85",x"E7", -- 0x1970
    x"8D",x"05",x"01",x"18",x"69",x"34",x"A2",x"1C", -- 0x1978
    x"A0",x"38",x"20",x"C2",x"AE",x"20",x"59",x"AB", -- 0x1980
    x"20",x"E5",x"A9",x"F0",x"A2",x"20",x"08",x"AA", -- 0x1988
    x"AD",x"04",x"01",x"85",x"EA",x"85",x"EB",x"A9", -- 0x1990
    x"02",x"85",x"E8",x"85",x"E9",x"AE",x"05",x"01", -- 0x1998
    x"BD",x"8D",x"AB",x"85",x"E9",x"A9",x"00",x"85", -- 0x19A0
    x"E7",x"20",x"59",x"AB",x"20",x"A1",x"AE",x"A2", -- 0x19A8
    x"FF",x"9A",x"4C",x"E3",x"A0",x"A0",x"05",x"A9", -- 0x19B0
    x"F0",x"20",x"95",x"AE",x"88",x"B9",x"C6",x"A9", -- 0x19B8
    x"8D",x"0C",x"90",x"D0",x"F2",x"60",x"00",x"E3", -- 0x19C0
    x"DB",x"D6",x"D2",x"C9",x"A2",x"06",x"86",x"21", -- 0x19C8
    x"BD",x"9B",x"AB",x"48",x"BC",x"95",x"AB",x"BD", -- 0x19D0
    x"8F",x"AB",x"AA",x"68",x"20",x"4F",x"AE",x"A6", -- 0x19D8
    x"21",x"CA",x"10",x"EA",x"60",x"A9",x"EF",x"20", -- 0x19E0
    x"EB",x"AC",x"29",x"80",x"D0",x"17",x"F0",x"09", -- 0x19E8
    x"A9",x"BF",x"20",x"EB",x"AC",x"29",x"80",x"D0", -- 0x19F0
    x"0C",x"A9",x"01",x"60",x"A9",x"DF",x"20",x"EB", -- 0x19F8
    x"AC",x"29",x"80",x"F0",x"F4",x"A9",x"00",x"60", -- 0x1A00
    x"20",x"93",x"AE",x"20",x"E5",x"A9",x"D0",x"F8", -- 0x1A08
    x"60",x"20",x"A1",x"AE",x"A9",x"2F",x"8D",x"0E", -- 0x1A10
    x"90",x"A6",x"E7",x"D6",x"E8",x"30",x"25",x"20", -- 0x1A18
    x"33",x"AB",x"20",x"D1",x"AB",x"A2",x"0A",x"20", -- 0x1A20
    x"93",x"AE",x"20",x"93",x"AE",x"8A",x"48",x"29", -- 0x1A28
    x"01",x"F0",x"06",x"20",x"B2",x"AB",x"4C",x"3C", -- 0x1A30
    x"AA",x"20",x"A1",x"AB",x"68",x"AA",x"CA",x"10", -- 0x1A38
    x"E6",x"4C",x"20",x"A1",x"20",x"D1",x"AB",x"A6", -- 0x1A40
    x"E7",x"A9",x"FF",x"95",x"E8",x"A0",x"08",x"84", -- 0x1A48
    x"0E",x"A2",x"18",x"86",x"0D",x"20",x"CD",x"AD", -- 0x1A50
    x"32",x"31",x"30",x"2E",x"16",x"16",x"2D",x"2C", -- 0x1A58
    x"2E",x"2A",x"00",x"20",x"A1",x"AE",x"A9",x"32", -- 0x1A60
    x"85",x"00",x"20",x"33",x"AB",x"A2",x"0A",x"20", -- 0x1A68
    x"93",x"AE",x"CA",x"D0",x"FA",x"A2",x"18",x"86", -- 0x1A70
    x"0D",x"A0",x"08",x"84",x"0E",x"20",x"CD",x"AD", -- 0x1A78
    x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16", -- 0x1A80
    x"16",x"16",x"00",x"4C",x"22",x"AA",x"A0",x"02", -- 0x1A88
    x"A9",x"00",x"19",x"EE",x"00",x"19",x"F0",x"00", -- 0x1A90
    x"19",x"F4",x"00",x"88",x"10",x"F4",x"24",x"E8", -- 0x1A98
    x"D0",x"03",x"20",x"66",x"B0",x"A0",x"01",x"84", -- 0x1AA0
    x"0C",x"E6",x"0C",x"A5",x"0C",x"C9",x"14",x"F0", -- 0x1AA8
    x"23",x"0A",x"0A",x"0A",x"A8",x"A2",x"00",x"20", -- 0x1AB0
    x"CD",x"AD",x"16",x"16",x"16",x"16",x"16",x"16", -- 0x1AB8
    x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16", -- 0x1AC0
    x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16", -- 0x1AC8
    x"00",x"4C",x"A9",x"AA",x"A2",x"02",x"A0",x"04", -- 0x1AD0
    x"A9",x"07",x"20",x"4F",x"AE",x"20",x"59",x"AB", -- 0x1AD8
    x"A2",x"10",x"A0",x"28",x"20",x"CD",x"AD",x"1B", -- 0x1AE0
    x"34",x"26",x"24",x"22",x"31",x"2A",x"22",x"16", -- 0x1AE8
    x"32",x"31",x"30",x"2E",x"00",x"A2",x"10",x"A0", -- 0x1AF0
    x"40",x"20",x"CD",x"AD",x"1B",x"38",x"26",x"2D", -- 0x1AF8
    x"28",x"22",x"20",x"2D",x"29",x"24",x"00",x"20", -- 0x1B00
    x"70",x"AB",x"20",x"22",x"AE",x"A5",x"0C",x"F0", -- 0x1B08
    x"10",x"20",x"E5",x"A9",x"D0",x"0B",x"20",x"F0", -- 0x1B10
    x"A9",x"F0",x"EC",x"20",x"59",x"AB",x"4C",x"71", -- 0x1B18
    x"A8",x"20",x"59",x"AB",x"20",x"90",x"A9",x"A2", -- 0x1B20
    x"FF",x"9A",x"4C",x"E3",x"A0",x"A2",x"FF",x"9A", -- 0x1B28
    x"4C",x"44",x"A0",x"A5",x"E7",x"49",x"01",x"AA", -- 0x1B30
    x"B5",x"E8",x"30",x"14",x"86",x"E7",x"A2",x"1D", -- 0x1B38
    x"B5",x"C9",x"A8",x"BD",x"E1",x"1F",x"95",x"C9", -- 0x1B40
    x"98",x"9D",x"E1",x"1F",x"CA",x"10",x"F1",x"60", -- 0x1B48
    x"A6",x"E7",x"B5",x"E8",x"10",x"36",x"4C",x"8E", -- 0x1B50
    x"AA",x"A9",x"0E",x"8D",x"0F",x"90",x"A9",x"2F", -- 0x1B58
    x"8D",x"0E",x"90",x"A9",x"00",x"85",x"A9",x"85", -- 0x1B60
    x"9E",x"85",x"9F",x"A9",x"24",x"85",x"A0",x"60", -- 0x1B68
    x"E6",x"9E",x"D0",x"18",x"E6",x"9F",x"D0",x"14", -- 0x1B70
    x"A5",x"A9",x"D0",x"04",x"C6",x"A0",x"D0",x"0C", -- 0x1B78
    x"A2",x"07",x"86",x"A9",x"20",x"FF",x"AD",x"09", -- 0x1B80
    x"08",x"8D",x"0F",x"90",x"60",x"FF",x"02",x"00", -- 0x1B88
    x"01",x"02",x"07",x"08",x"0A",x"00",x"01",x"06", -- 0x1B90
    x"07",x"09",x"0A",x"07",x"06",x"07",x"0F",x"03", -- 0x1B98
    x"07",x"A2",x"38",x"A0",x"A8",x"20",x"CD",x"AD", -- 0x1BA0
    x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16", -- 0x1BA8
    x"00",x"60",x"A2",x"38",x"A0",x"A8",x"20",x"CD", -- 0x1BB0
    x"AD",x"28",x"27",x"31",x"19",x"2E",x"2A",x"00", -- 0x1BB8
    x"A2",x"54",x"A0",x"A8",x"A5",x"E7",x"18",x"69", -- 0x1BC0
    x"34",x"20",x"C2",x"AE",x"60",x"A6",x"E7",x"F6", -- 0x1BC8
    x"E8",x"20",x"B2",x"AB",x"A2",x"00",x"A0",x"A8", -- 0x1BD0
    x"20",x"CD",x"AD",x"16",x"16",x"16",x"16",x"16", -- 0x1BD8
    x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16", -- 0x1BE0
    x"16",x"00",x"A0",x"A8",x"84",x"0E",x"A2",x"00", -- 0x1BE8
    x"86",x"0D",x"A4",x"E7",x"B6",x"E8",x"86",x"A3", -- 0x1BF0
    x"30",x"2E",x"F0",x"16",x"C6",x"A3",x"E0",x"0D", -- 0x1BF8
    x"90",x"04",x"A2",x"0C",x"86",x"A3",x"A9",x"15", -- 0x1C00
    x"20",x"C6",x"AE",x"A5",x"0D",x"18",x"69",x"04", -- 0x1C08
    x"85",x"0D",x"A9",x"16",x"20",x"C6",x"AE",x"C6", -- 0x1C10
    x"A3",x"10",x"EB",x"A6",x"E7",x"B5",x"E8",x"C9", -- 0x1C18
    x"0D",x"90",x"05",x"A9",x"25",x"4C",x"C6",x"AE", -- 0x1C20
    x"60",x"20",x"A1",x"AE",x"A6",x"E7",x"A5",x"6C", -- 0x1C28
    x"C9",x"08",x"F0",x"02",x"F6",x"6C",x"F8",x"B5", -- 0x1C30
    x"EA",x"18",x"69",x"01",x"95",x"EA",x"D8",x"20", -- 0x1C38
    x"48",x"AC",x"A2",x"FF",x"9A",x"4C",x"F8",x"A0", -- 0x1C40
    x"A9",x"A0",x"85",x"0E",x"A9",x"58",x"85",x"0D", -- 0x1C48
    x"A9",x"16",x"20",x"C6",x"AE",x"A5",x"0D",x"38", -- 0x1C50
    x"E9",x"04",x"10",x"F2",x"A2",x"54",x"86",x"0D", -- 0x1C58
    x"A6",x"E7",x"B5",x"EA",x"F8",x"18",x"69",x"01", -- 0x1C60
    x"D8",x"4A",x"4A",x"4A",x"4A",x"F0",x"12",x"85", -- 0x1C68
    x"21",x"A9",x"17",x"20",x"C6",x"AE",x"A5",x"0D", -- 0x1C70
    x"38",x"E9",x"04",x"85",x"0D",x"C6",x"21",x"D0", -- 0x1C78
    x"F0",x"A6",x"E7",x"B5",x"EA",x"F8",x"18",x"69", -- 0x1C80
    x"01",x"D8",x"29",x"0F",x"F0",x"12",x"85",x"21", -- 0x1C88
    x"A9",x"18",x"20",x"C6",x"AE",x"A5",x"0D",x"38", -- 0x1C90
    x"E9",x"04",x"85",x"0D",x"C6",x"21",x"D0",x"F0", -- 0x1C98
    x"60",x"20",x"F0",x"A9",x"F0",x"03",x"4C",x"71", -- 0x1CA0
    x"A8",x"20",x"E5",x"A9",x"F0",x"09",x"20",x"90", -- 0x1CA8
    x"A9",x"A2",x"FF",x"9A",x"4C",x"E3",x"A0",x"20", -- 0x1CB0
    x"DE",x"AC",x"90",x"3A",x"A9",x"20",x"8D",x"0E", -- 0x1CB8
    x"90",x"20",x"93",x"AE",x"20",x"D8",x"AC",x"20", -- 0x1CC0
    x"70",x"AB",x"20",x"DE",x"AC",x"90",x"F8",x"20", -- 0x1CC8
    x"D8",x"AC",x"20",x"93",x"AE",x"4C",x"59",x"AB", -- 0x1CD0
    x"20",x"DE",x"AC",x"B0",x"FB",x"60",x"A9",x"EF", -- 0x1CD8
    x"20",x"EB",x"AC",x"29",x"01",x"D0",x"02",x"38", -- 0x1CE0
    x"60",x"18",x"60",x"8D",x"20",x"91",x"AD",x"21", -- 0x1CE8
    x"91",x"CD",x"21",x"91",x"D0",x"F8",x"60",x"48", -- 0x1CF0
    x"86",x"00",x"A5",x"E7",x"0A",x"18",x"65",x"E7", -- 0x1CF8
    x"AA",x"68",x"F8",x"18",x"75",x"EE",x"95",x"EE", -- 0x1D00
    x"A5",x"00",x"75",x"EF",x"95",x"EF",x"A9",x"00", -- 0x1D08
    x"75",x"F0",x"95",x"F0",x"D8",x"86",x"0C",x"A4", -- 0x1D10
    x"E7",x"B5",x"EF",x"C9",x"70",x"90",x"0E",x"B9", -- 0x1D18
    x"EC",x"00",x"D0",x"07",x"A6",x"E7",x"F6",x"EC", -- 0x1D20
    x"20",x"CD",x"AB",x"A6",x"0C",x"E8",x"E8",x"86", -- 0x1D28
    x"00",x"A0",x"02",x"B5",x"EE",x"D9",x"F4",x"00", -- 0x1D30
    x"90",x"15",x"F0",x"02",x"B0",x"04",x"CA",x"88", -- 0x1D38
    x"10",x"F1",x"A6",x"00",x"A0",x"02",x"B5",x"EE", -- 0x1D40
    x"99",x"F4",x"00",x"CA",x"88",x"10",x"F7",x"A2", -- 0x1D48
    x"20",x"A0",x"00",x"A9",x"F4",x"85",x"22",x"A9", -- 0x1D50
    x"00",x"85",x"23",x"A9",x"02",x"20",x"80",x"AD", -- 0x1D58
    x"A9",x"EE",x"85",x"22",x"A9",x"00",x"85",x"23", -- 0x1D60
    x"A2",x"00",x"A0",x"00",x"A9",x"02",x"20",x"80", -- 0x1D68
    x"AD",x"AD",x"05",x"01",x"F0",x"56",x"A9",x"F1", -- 0x1D70
    x"85",x"22",x"A2",x"40",x"A0",x"00",x"A9",x"02", -- 0x1D78
    x"86",x"0D",x"84",x"0E",x"85",x"24",x"A2",x"00", -- 0x1D80
    x"86",x"AA",x"A4",x"24",x"B1",x"22",x"48",x"4A", -- 0x1D88
    x"4A",x"4A",x"4A",x"18",x"69",x"33",x"C9",x"33", -- 0x1D90
    x"D0",x"04",x"A6",x"AA",x"F0",x"07",x"A2",x"01", -- 0x1D98
    x"86",x"AA",x"20",x"C6",x"AE",x"A5",x"0D",x"18", -- 0x1DA0
    x"69",x"04",x"85",x"0D",x"68",x"29",x"0F",x"18", -- 0x1DA8
    x"69",x"33",x"C9",x"33",x"D0",x"04",x"A6",x"AA", -- 0x1DB0
    x"F0",x"07",x"A2",x"01",x"86",x"AA",x"20",x"C6", -- 0x1DB8
    x"AE",x"A5",x"0D",x"18",x"69",x"04",x"85",x"0D", -- 0x1DC0
    x"C6",x"24",x"10",x"BE",x"60",x"86",x"0D",x"84", -- 0x1DC8
    x"0E",x"68",x"85",x"2C",x"68",x"85",x"2D",x"D0", -- 0x1DD0
    x"10",x"A0",x"00",x"B1",x"2C",x"F0",x"12",x"20", -- 0x1DD8
    x"C6",x"AE",x"A5",x"0D",x"18",x"69",x"04",x"85", -- 0x1DE0
    x"0D",x"E6",x"2C",x"D0",x"EC",x"E6",x"2D",x"D0", -- 0x1DE8
    x"E8",x"A5",x"2D",x"48",x"A5",x"2C",x"48",x"60", -- 0x1DF0
    x"A5",x"0C",x"29",x"10",x"D0",x"FA",x"60",x"AD", -- 0x1DF8
    x"04",x"90",x"6D",x"01",x"01",x"EE",x"03",x"01", -- 0x1E00
    x"EE",x"00",x"01",x"AC",x"03",x"01",x"71",x"FF", -- 0x1E08
    x"6D",x"04",x"90",x"8D",x"01",x"01",x"3D",x"1A", -- 0x1E10
    x"AE",x"60",x"01",x"03",x"07",x"0F",x"1F",x"3F", -- 0x1E18
    x"7F",x"FF",x"A0",x"03",x"A9",x"FF",x"C0",x"02", -- 0x1E20
    x"F0",x"09",x"8D",x"22",x"91",x"AD",x"11",x"91", -- 0x1E28
    x"4C",x"3A",x"AE",x"4A",x"8D",x"22",x"91",x"AD", -- 0x1E30
    x"20",x"91",x"39",x"4B",x"AE",x"99",x"08",x"00", -- 0x1E38
    x"88",x"10",x"E1",x"AD",x"11",x"91",x"29",x"20", -- 0x1E40
    x"85",x"0C",x"60",x"10",x"04",x"80",x"08",x"86", -- 0x1E48
    x"06",x"84",x"07",x"48",x"20",x"8A",x"AE",x"A0", -- 0x1E50
    x"15",x"68",x"91",x"04",x"88",x"10",x"FB",x"A4", -- 0x1E58
    x"07",x"C4",x"06",x"F0",x"24",x"88",x"10",x"E9", -- 0x1E60
    x"A9",x"10",x"85",x"03",x"A9",x"00",x"85",x"02", -- 0x1E68
    x"A8",x"A2",x"0F",x"91",x"02",x"99",x"20",x"1E", -- 0x1E70
    x"C8",x"D0",x"F8",x"E6",x"03",x"CA",x"D0",x"F3", -- 0x1E78
    x"60",x"B1",x"F7",x"85",x"02",x"B1",x"F9",x"85", -- 0x1E80
    x"03",x"60",x"B1",x"FB",x"85",x"04",x"B1",x"FD", -- 0x1E88
    x"85",x"05",x"60",x"A9",x"FF",x"38",x"48",x"E9", -- 0x1E90
    x"01",x"D0",x"FC",x"68",x"E9",x"01",x"D0",x"F6", -- 0x1E98
    x"60",x"20",x"B0",x"AE",x"20",x"B6",x"AE",x"20", -- 0x1EA0
    x"BC",x"AE",x"A9",x"00",x"8D",x"0D",x"90",x"60", -- 0x1EA8
    x"A9",x"00",x"8D",x"0A",x"90",x"60",x"A9",x"00", -- 0x1EB0
    x"8D",x"0B",x"90",x"60",x"A9",x"00",x"8D",x"0C", -- 0x1EB8
    x"90",x"60",x"86",x"0D",x"84",x"0E",x"A6",x"0D", -- 0x1EC0
    x"85",x"18",x"8A",x"29",x"03",x"85",x"19",x"8A", -- 0x1EC8
    x"4A",x"4A",x"85",x"14",x"A5",x"18",x"0A",x"A8", -- 0x1ED0
    x"B9",x"E4",x"B1",x"85",x"1A",x"C8",x"B9",x"E4", -- 0x1ED8
    x"B1",x"85",x"1B",x"A0",x"00",x"B1",x"1A",x"85", -- 0x1EE0
    x"11",x"C8",x"B1",x"1A",x"85",x"12",x"A5",x"1A", -- 0x1EE8
    x"18",x"69",x"02",x"85",x"15",x"A5",x"1B",x"69", -- 0x1EF0
    x"00",x"85",x"16",x"A9",x"00",x"85",x"1C",x"A5", -- 0x1EF8
    x"12",x"85",x"17",x"A5",x"0E",x"85",x"1D",x"A4", -- 0x1F00
    x"14",x"C0",x"16",x"B0",x"4A",x"20",x"81",x"AE", -- 0x1F08
    x"A5",x"17",x"C5",x"12",x"F0",x"42",x"C9",x"01", -- 0x1F10
    x"F0",x"42",x"A2",x"04",x"A4",x"11",x"84",x"13", -- 0x1F18
    x"A9",x"00",x"A4",x"1C",x"20",x"6D",x"AF",x"A4", -- 0x1F20
    x"1D",x"48",x"AD",x"02",x"01",x"F0",x"08",x"10", -- 0x1F28
    x"0C",x"68",x"31",x"02",x"4C",x"47",x"AF",x"68", -- 0x1F30
    x"11",x"02",x"4C",x"47",x"AF",x"B1",x"02",x"3D", -- 0x1F38
    x"64",x"AF",x"85",x"00",x"68",x"05",x"00",x"91", -- 0x1F40
    x"02",x"E6",x"1C",x"E6",x"1D",x"C6",x"13",x"D0", -- 0x1F48
    x"CF",x"E6",x"14",x"C6",x"17",x"D0",x"AC",x"60", -- 0x1F50
    x"A6",x"19",x"10",x"C0",x"A9",x"05",x"18",x"65", -- 0x1F58
    x"19",x"AA",x"D0",x"B8",x"00",x"C0",x"F0",x"FC", -- 0x1F60
    x"00",x"FF",x"3F",x"0F",x"03",x"85",x"0F",x"86", -- 0x1F68
    x"10",x"E0",x"04",x"90",x"1B",x"F0",x"21",x"98", -- 0x1F70
    x"38",x"E5",x"11",x"A8",x"B1",x"15",x"A8",x"A5", -- 0x1F78
    x"19",x"18",x"69",x"FC",x"AA",x"98",x"0A",x"0A", -- 0x1F80
    x"E8",x"D0",x"FB",x"05",x"0F",x"A6",x"10",x"60", -- 0x1F88
    x"B1",x"15",x"20",x"A4",x"AF",x"4C",x"8B",x"AF", -- 0x1F90
    x"B1",x"15",x"20",x"A4",x"AF",x"05",x"0F",x"85", -- 0x1F98
    x"0F",x"4C",x"77",x"AF",x"A6",x"19",x"F0",x"05", -- 0x1FA0
    x"4A",x"4A",x"CA",x"D0",x"FB",x"60",x"00",x"0A", -- 0x1FA8
    x"0C",x"0F",x"0E",x"0D",x"0E",x"0D",x"0C",x"0D", -- 0x1FB0
    x"0C",x"0B",x"00",x"00",x"00",x"01",x"01",x"02", -- 0x1FB8
    x"02",x"07",x"00",x"00",x"90",x"40",x"40",x"40", -- 0x1FC0
    x"40",x"40",x"00",x"1A",x"19",x"1B",x"00",x"17", -- 0x1FC8
    x"18",x"16",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FD0
    x"20",x"20",x"31",x"39",x"38",x"34",x"20",x"20", -- 0x1FD8
    x"44",x"45",x"53",x"49",x"47",x"4E",x"45",x"52", -- 0x1FE0
    x"53",x"4F",x"46",x"54",x"57",x"41",x"52",x"45", -- 0x1FE8
    x"42",x"49",x"4C",x"4C",x"20",x"42",x"4F",x"47", -- 0x1FF0
    x"45",x"4E",x"52",x"45",x"49",x"46",x"20",x"36"  -- 0x1FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
