-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity cart_rom is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of cart_rom is


  type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"12",x"A0",x"09",x"A0",x"41",x"30",x"C3",x"C2", -- 0x0000
    x"CD",x"D8",x"68",x"A8",x"68",x"AA",x"68",x"4C", -- 0x0008
    x"35",x"A0",x"20",x"8D",x"FD",x"20",x"F9",x"FD", -- 0x0010
    x"20",x"18",x"E5",x"20",x"8A",x"FF",x"AD",x"01", -- 0x0018
    x"90",x"E9",x"04",x"8D",x"01",x"90",x"A9",x"95", -- 0x0020
    x"8D",x"02",x"90",x"A9",x"B0",x"8D",x"03",x"90", -- 0x0028
    x"A2",x"FF",x"8E",x"05",x"90",x"78",x"A2",x"09", -- 0x0030
    x"A0",x"AA",x"8E",x"14",x"03",x"8C",x"15",x"03", -- 0x0038
    x"58",x"A9",x"00",x"85",x"FC",x"A9",x"AC",x"85", -- 0x0040
    x"FD",x"A9",x"00",x"85",x"FE",x"A9",x"1A",x"85", -- 0x0048
    x"FF",x"A0",x"00",x"B1",x"FC",x"91",x"FE",x"C8", -- 0x0050
    x"D0",x"F9",x"E6",x"FD",x"E6",x"FF",x"A5",x"FF", -- 0x0058
    x"C9",x"1E",x"D0",x"EF",x"98",x"99",x"0A",x"90", -- 0x0060
    x"C8",x"C0",x"04",x"D0",x"F8",x"A9",x"8F",x"8D", -- 0x0068
    x"0E",x"90",x"20",x"06",x"A7",x"A2",x"15",x"BD", -- 0x0070
    x"E3",x"AD",x"9D",x"E3",x"1F",x"A9",x"03",x"9D", -- 0x0078
    x"E3",x"97",x"CA",x"10",x"F2",x"A9",x"09",x"8D", -- 0x0080
    x"F1",x"97",x"8D",x"F2",x"97",x"20",x"EC",x"A6", -- 0x0088
    x"A0",x"00",x"84",x"45",x"20",x"AA",x"AB",x"A0", -- 0x0090
    x"0A",x"8C",x"A1",x"02",x"A5",x"44",x"29",x"7F", -- 0x0098
    x"D0",x"30",x"AE",x"0F",x"90",x"E8",x"8A",x"29", -- 0x00A0
    x"07",x"AA",x"09",x"08",x"8D",x"0F",x"90",x"20", -- 0x00A8
    x"81",x"A7",x"E6",x"49",x"A6",x"49",x"E0",x"0D", -- 0x00B0
    x"90",x"06",x"86",x"3B",x"A2",x"00",x"86",x"49", -- 0x00B8
    x"BD",x"55",x"AE",x"8D",x"1B",x"1F",x"BD",x"62", -- 0x00C0
    x"AE",x"8D",x"1B",x"97",x"A9",x"40",x"85",x"39", -- 0x00C8
    x"85",x"3A",x"A6",x"A2",x"E8",x"E8",x"E4",x"A2", -- 0x00D0
    x"D0",x"FC",x"AD",x"A1",x"02",x"49",x"1E",x"8D", -- 0x00D8
    x"A1",x"02",x"20",x"FD",x"A2",x"20",x"15",x"A8", -- 0x00E0
    x"20",x"E4",x"FF",x"C9",x"85",x"F0",x"0C",x"A9", -- 0x00E8
    x"FF",x"8D",x"22",x"91",x"AD",x"11",x"91",x"29", -- 0x00F0
    x"20",x"D0",x"A1",x"A9",x"09",x"85",x"3C",x"A9", -- 0x00F8
    x"03",x"85",x"45",x"A0",x"FF",x"84",x"49",x"20", -- 0x0100
    x"AA",x"AB",x"A2",x"00",x"86",x"47",x"A9",x"B0", -- 0x0108
    x"9D",x"06",x"1A",x"E8",x"E0",x"06",x"D0",x"F6", -- 0x0110
    x"20",x"06",x"A7",x"20",x"EC",x"A6",x"A9",x"1C", -- 0x0118
    x"8D",x"C2",x"02",x"A9",x"A8",x"8D",x"BA",x"02", -- 0x0120
    x"A9",x"1F",x"8D",x"A1",x"02",x"A2",x"0C",x"A9", -- 0x0128
    x"08",x"20",x"99",x"AB",x"CA",x"10",x"F8",x"A2", -- 0x0130
    x"05",x"BD",x"77",x"C3",x"29",x"BF",x"09",x"80", -- 0x0138
    x"9D",x"18",x"1F",x"A9",x"07",x"9D",x"18",x"97", -- 0x0140
    x"A9",x"98",x"9D",x"BA",x"02",x"CA",x"D0",x"E9", -- 0x0148
    x"A9",x"C8",x"8D",x"BA",x"02",x"A2",x"18",x"A9", -- 0x0150
    x"08",x"20",x"99",x"AB",x"CA",x"10",x"F8",x"A2", -- 0x0158
    x"00",x"A9",x"20",x"9D",x"19",x"1F",x"E8",x"E0", -- 0x0160
    x"05",x"D0",x"F8",x"A2",x"00",x"86",x"3A",x"86", -- 0x0168
    x"3B",x"86",x"3D",x"A2",x"02",x"86",x"43",x"86", -- 0x0170
    x"42",x"AD",x"8D",x"02",x"D0",x"FB",x"AD",x"1B", -- 0x0178
    x"1F",x"C9",x"21",x"90",x"08",x"A6",x"49",x"BD", -- 0x0180
    x"62",x"AE",x"8D",x"1B",x"97",x"A9",x"0C",x"38", -- 0x0188
    x"E5",x"49",x"90",x"04",x"C9",x"03",x"B0",x"02", -- 0x0190
    x"A9",x"03",x"A8",x"E8",x"D0",x"FD",x"88",x"D0", -- 0x0198
    x"FA",x"84",x"00",x"84",x"01",x"A5",x"43",x"85", -- 0x01A0
    x"40",x"A6",x"42",x"8C",x"13",x"91",x"A9",x"7F", -- 0x01A8
    x"8D",x"22",x"91",x"AD",x"20",x"91",x"29",x"80", -- 0x01B0
    x"D0",x"02",x"A2",x"00",x"A9",x"FF",x"8D",x"22", -- 0x01B8
    x"91",x"AC",x"11",x"91",x"98",x"29",x"08",x"D0", -- 0x01C0
    x"02",x"A2",x"01",x"98",x"29",x"10",x"D0",x"02", -- 0x01C8
    x"A2",x"02",x"98",x"29",x"04",x"D0",x"02",x"A2", -- 0x01D0
    x"03",x"86",x"42",x"8A",x"85",x"41",x"20",x"A7", -- 0x01D8
    x"A7",x"B0",x"07",x"A5",x"42",x"85",x"43",x"18", -- 0x01E0
    x"90",x"07",x"A5",x"43",x"85",x"41",x"20",x"A7", -- 0x01E8
    x"A7",x"AD",x"A2",x"02",x"D0",x"05",x"A9",x"9E", -- 0x01F0
    x"8D",x"A2",x"02",x"C9",x"A0",x"D0",x"05",x"A9", -- 0x01F8
    x"00",x"8D",x"A2",x"02",x"A2",x"B0",x"AD",x"A2", -- 0x0200
    x"02",x"0D",x"A3",x"02",x"29",x"02",x"D0",x"09", -- 0x0208
    x"A5",x"43",x"0A",x"0A",x"0A",x"18",x"69",x"B8", -- 0x0210
    x"AA",x"8E",x"BA",x"02",x"A2",x"00",x"AD",x"A2", -- 0x0218
    x"02",x"29",x"07",x"C9",x"04",x"D0",x"0B",x"E8", -- 0x0220
    x"A5",x"43",x"49",x"02",x"A8",x"F0",x"15",x"88", -- 0x0228
    x"D0",x"12",x"AD",x"A3",x"02",x"29",x"07",x"C9", -- 0x0230
    x"03",x"D0",x"09",x"E8",x"A4",x"43",x"C0",x"01", -- 0x0238
    x"F0",x"02",x"A0",x"00",x"E0",x"00",x"D0",x"03", -- 0x0240
    x"4C",x"ED",x"A2",x"B9",x"DD",x"02",x"C9",x"20", -- 0x0248
    x"D0",x"03",x"4C",x"79",x"A1",x"AA",x"A9",x"20", -- 0x0250
    x"99",x"DD",x"02",x"E0",x"1E",x"D0",x"0A",x"A9", -- 0x0258
    x"01",x"85",x"3F",x"85",x"3D",x"A9",x"0A",x"85", -- 0x0260
    x"3E",x"E0",x"21",x"90",x"17",x"E0",x"29",x"B0", -- 0x0268
    x"7C",x"8A",x"38",x"E9",x"21",x"AA",x"BD",x"F8", -- 0x0270
    x"AD",x"85",x"3F",x"A9",x"09",x"85",x"3E",x"85", -- 0x0278
    x"3C",x"18",x"90",x"69",x"E0",x"1F",x"D0",x"0C", -- 0x0280
    x"A9",x"05",x"85",x"3F",x"A9",x"0A",x"85",x"3E", -- 0x0288
    x"85",x"3B",x"F0",x"59",x"E6",x"4A",x"A5",x"4A", -- 0x0290
    x"C9",x"AA",x"D0",x"51",x"A9",x"A8",x"8D",x"BA", -- 0x0298
    x"02",x"A9",x"80",x"20",x"99",x"AB",x"A9",x"00", -- 0x02A0
    x"85",x"44",x"C6",x"44",x"A5",x"44",x"29",x"07", -- 0x02A8
    x"AA",x"20",x"81",x"A7",x"A5",x"44",x"29",x"1F", -- 0x02B0
    x"D0",x"08",x"AD",x"A1",x"02",x"49",x"1E",x"8D", -- 0x02B8
    x"A1",x"02",x"A2",x"04",x"A9",x"70",x"9D",x"BA", -- 0x02C0
    x"02",x"CA",x"D0",x"FA",x"20",x"15",x"A8",x"A5", -- 0x02C8
    x"44",x"C9",x"06",x"D0",x"D5",x"A9",x"40",x"20", -- 0x02D0
    x"99",x"AB",x"A2",x"03",x"B5",x"4B",x"A4",x"49", -- 0x02D8
    x"C8",x"4A",x"88",x"D0",x"FC",x"95",x"4B",x"CA", -- 0x02E0
    x"10",x"F2",x"4C",x"18",x"A1",x"20",x"E4",x"FF", -- 0x02E8
    x"C9",x"03",x"F0",x"A8",x"20",x"FD",x"A2",x"20", -- 0x02F0
    x"15",x"A8",x"4C",x"79",x"A1",x"A5",x"3A",x"D0", -- 0x02F8
    x"24",x"A5",x"4A",x"C9",x"4B",x"F0",x"04",x"C9", -- 0x0300
    x"7D",x"D0",x"1A",x"A6",x"49",x"E0",x"0C",x"90", -- 0x0308
    x"02",x"A2",x"0C",x"BD",x"55",x"AE",x"8D",x"1B", -- 0x0310
    x"1F",x"BD",x"62",x"AE",x"8D",x"1B",x"97",x"A9", -- 0x0318
    x"FA",x"85",x"39",x"85",x"3A",x"A5",x"39",x"F0", -- 0x0320
    x"09",x"C6",x"39",x"D0",x"05",x"A9",x"20",x"8D", -- 0x0328
    x"1B",x"1F",x"A5",x"4A",x"C9",x"4C",x"F0",x"04", -- 0x0330
    x"C9",x"7E",x"D0",x"04",x"A9",x"00",x"85",x"3A", -- 0x0338
    x"A5",x"3B",x"F0",x"3C",x"A9",x"00",x"85",x"3B", -- 0x0340
    x"A9",x"02",x"85",x"70",x"A6",x"49",x"8A",x"29", -- 0x0348
    x"07",x"F0",x"05",x"E0",x"10",x"B0",x"0C",x"8A", -- 0x0350
    x"0A",x"0A",x"29",x"3F",x"49",x"3F",x"E0",x"05", -- 0x0358
    x"90",x"01",x"4A",x"85",x"10",x"A0",x"04",x"B6", -- 0x0360
    x"4A",x"D0",x"12",x"A9",x"06",x"99",x"B2",x"02", -- 0x0368
    x"A9",x"A0",x"99",x"BA",x"02",x"B9",x"4E",x"00", -- 0x0370
    x"49",x"02",x"99",x"4E",x"00",x"88",x"D0",x"E7", -- 0x0378
    x"A0",x"08",x"A5",x"45",x"F0",x"32",x"AD",x"A2", -- 0x0380
    x"02",x"D9",x"A2",x"02",x"D0",x"13",x"AD",x"A3", -- 0x0388
    x"02",x"38",x"F9",x"A3",x"02",x"B0",x"02",x"49", -- 0x0390
    x"FF",x"C9",x"05",x"B0",x"04",x"A2",x"FF",x"D0", -- 0x0398
    x"1E",x"AD",x"A3",x"02",x"D9",x"A3",x"02",x"D0", -- 0x03A0
    x"0F",x"AD",x"A2",x"02",x"38",x"F9",x"A2",x"02", -- 0x03A8
    x"B0",x"02",x"49",x"FF",x"C9",x"05",x"90",x"07", -- 0x03B0
    x"88",x"88",x"D0",x"C6",x"4C",x"FC",x"A4",x"98", -- 0x03B8
    x"4A",x"AA",x"BD",x"BA",x"02",x"C9",x"70",x"F0", -- 0x03C0
    x"EF",x"C9",x"A0",x"D0",x"64",x"A9",x"09",x"85", -- 0x03C8
    x"3E",x"A5",x"70",x"85",x"3F",x"0A",x"85",x"70", -- 0x03D0
    x"98",x"48",x"8A",x"48",x"A9",x"D0",x"8D",x"0A", -- 0x03D8
    x"90",x"AD",x"A1",x"02",x"5D",x"FB",x"AB",x"8D", -- 0x03E0
    x"A1",x"02",x"A6",x"10",x"A9",x"01",x"20",x"99", -- 0x03E8
    x"AB",x"A9",x"A8",x"8D",x"BA",x"02",x"A9",x"01", -- 0x03F0
    x"20",x"99",x"AB",x"A5",x"A2",x"18",x"69",x"20", -- 0x03F8
    x"A4",x"A2",x"C8",x"C4",x"A2",x"D0",x"FC",x"86", -- 0x0400
    x"10",x"EE",x"0A",x"90",x"C5",x"A2",x"D0",x"F0", -- 0x0408
    x"A9",x"00",x"8D",x"0A",x"90",x"68",x"AA",x"68", -- 0x0410
    x"A8",x"A9",x"70",x"9D",x"BA",x"02",x"AD",x"A1", -- 0x0418
    x"02",x"5D",x"FB",x"AB",x"8D",x"A1",x"02",x"CA", -- 0x0420
    x"BD",x"51",x"AE",x"9D",x"B3",x"02",x"4C",x"B8", -- 0x0428
    x"A3",x"68",x"68",x"A2",x"06",x"A9",x"10",x"20", -- 0x0430
    x"99",x"AB",x"CA",x"10",x"F8",x"A9",x"01",x"8D", -- 0x0438
    x"A1",x"02",x"A9",x"B0",x"8D",x"BA",x"02",x"A2", -- 0x0440
    x"01",x"BD",x"50",x"AE",x"9D",x"B2",x"02",x"A9", -- 0x0448
    x"80",x"9D",x"BA",x"02",x"E8",x"E0",x"05",x"D0", -- 0x0450
    x"F0",x"A9",x"F0",x"8D",x"0C",x"90",x"A9",x"20", -- 0x0458
    x"85",x"44",x"AD",x"BA",x"02",x"C9",x"D0",x"90", -- 0x0460
    x"05",x"EE",x"0C",x"90",x"A9",x"B0",x"18",x"69", -- 0x0468
    x"08",x"8D",x"BA",x"02",x"CE",x"0C",x"90",x"CE", -- 0x0470
    x"0C",x"90",x"CE",x"0C",x"90",x"A9",x"04",x"20", -- 0x0478
    x"99",x"AB",x"C6",x"44",x"D0",x"DC",x"A2",x"D8", -- 0x0480
    x"8E",x"BA",x"02",x"A9",x"0A",x"20",x"99",x"AB", -- 0x0488
    x"A2",x"E0",x"8E",x"BA",x"02",x"A9",x"08",x"20", -- 0x0490
    x"99",x"AB",x"A2",x"E8",x"8E",x"BA",x"02",x"A9", -- 0x0498
    x"06",x"20",x"99",x"AB",x"A9",x"00",x"8D",x"A1", -- 0x04A0
    x"02",x"8D",x"0C",x"90",x"A9",x"64",x"20",x"99", -- 0x04A8
    x"AB",x"C6",x"45",x"F0",x"37",x"A6",x"45",x"A9", -- 0x04B0
    x"1B",x"9D",x"E4",x"1F",x"A9",x"0A",x"20",x"99", -- 0x04B8
    x"AB",x"A9",x"1C",x"9D",x"E4",x"1F",x"A9",x"08", -- 0x04C0
    x"20",x"99",x"AB",x"A9",x"1D",x"9D",x"E4",x"1F", -- 0x04C8
    x"A9",x"01",x"8D",x"A1",x"02",x"A9",x"D8",x"8D", -- 0x04D0
    x"BA",x"02",x"20",x"EC",x"A6",x"A9",x"06",x"20", -- 0x04D8
    x"99",x"AB",x"A6",x"45",x"A9",x"20",x"9D",x"E4", -- 0x04E0
    x"1F",x"4C",x"1B",x"A1",x"A0",x"00",x"8C",x"A1", -- 0x04E8
    x"02",x"20",x"AA",x"AB",x"A9",x"F0",x"20",x"99", -- 0x04F0
    x"AB",x"4C",x"8D",x"A0",x"A9",x"04",x"85",x"00", -- 0x04F8
    x"A5",x"00",x"A8",x"0A",x"85",x"01",x"B6",x"4A", -- 0x0500
    x"F0",x"50",x"A5",x"44",x"29",x"03",x"F0",x"03", -- 0x0508
    x"CA",x"96",x"4A",x"A9",x"98",x"E0",x"10",x"90", -- 0x0510
    x"0B",x"8A",x"29",x"08",x"D0",x"04",x"A9",x"78", -- 0x0518
    x"D0",x"02",x"A9",x"88",x"99",x"BA",x"02",x"A6", -- 0x0520
    x"01",x"BD",x"A2",x"02",x"29",x"F8",x"9D",x"A2", -- 0x0528
    x"02",x"C6",x"00",x"D0",x"CB",x"E6",x"44",x"E6", -- 0x0530
    x"00",x"AD",x"A5",x"02",x"C9",x"58",x"F0",x"0D", -- 0x0538
    x"29",x"07",x"0D",x"A4",x"02",x"29",x"0F",x"F0", -- 0x0540
    x"B7",x"A5",x"3D",x"D0",x"01",x"60",x"A5",x"4A", -- 0x0548
    x"29",x"01",x"D0",x"F9",x"20",x"15",x"A8",x"4C", -- 0x0550
    x"FC",x"A4",x"B9",x"BA",x"02",x"C9",x"70",x"D0", -- 0x0558
    x"3D",x"A6",x"01",x"BD",x"A2",x"02",x"C9",x"50", -- 0x0560
    x"D0",x"0E",x"BD",x"A3",x"02",x"C9",x"48",x"D0", -- 0x0568
    x"07",x"FE",x"A3",x"02",x"A2",x"01",x"96",x"4E", -- 0x0570
    x"BD",x"A3",x"02",x"C9",x"58",x"D0",x"45",x"98", -- 0x0578
    x"0A",x"0A",x"0A",x"18",x"69",x"40",x"DD",x"A2", -- 0x0580
    x"02",x"D0",x"39",x"A9",x"98",x"99",x"BA",x"02", -- 0x0588
    x"B9",x"C3",x"AB",x"49",x"FF",x"4A",x"69",x"20", -- 0x0590
    x"99",x"4A",x"00",x"4C",x"31",x"A5",x"A5",x"44", -- 0x0598
    x"29",x"01",x"F0",x"07",x"B9",x"BA",x"02",x"C9", -- 0x05A0
    x"A0",x"F0",x"86",x"A6",x"01",x"BD",x"A2",x"02", -- 0x05A8
    x"C9",x"50",x"D0",x"10",x"BD",x"A3",x"02",x"C9", -- 0x05B0
    x"58",x"D0",x"09",x"DE",x"A3",x"02",x"A2",x"03", -- 0x05B8
    x"96",x"4E",x"D0",x"13",x"BD",x"A2",x"02",x"D0", -- 0x05C0
    x"04",x"A6",x"00",x"95",x"4E",x"C9",x"9F",x"D0", -- 0x05C8
    x"06",x"A6",x"00",x"A9",x"02",x"95",x"4E",x"A0", -- 0x05D0
    x"00",x"A2",x"04",x"96",x"60",x"C8",x"CA",x"D0", -- 0x05D8
    x"FA",x"A4",x"01",x"B9",x"A2",x"02",x"29",x"07", -- 0x05E0
    x"F0",x"07",x"B9",x"A3",x"02",x"29",x"07",x"D0", -- 0x05E8
    x"06",x"20",x"5A",x"A6",x"18",x"90",x"04",x"B6", -- 0x05F0
    x"4E",x"86",x"61",x"A0",x"00",x"84",x"04",x"B6", -- 0x05F8
    x"61",x"8A",x"A6",x"00",x"55",x"4E",x"C9",x"02", -- 0x0600
    x"F0",x"0F",x"B6",x"61",x"86",x"41",x"A4",x"00", -- 0x0608
    x"B6",x"4E",x"86",x"40",x"20",x"A7",x"A7",x"90", -- 0x0610
    x"14",x"E6",x"04",x"A4",x"04",x"C0",x"04",x"D0", -- 0x0618
    x"DE",x"A4",x"00",x"A5",x"40",x"49",x"02",x"99", -- 0x0620
    x"4E",x"00",x"4C",x"31",x"A5",x"A4",x"00",x"A6", -- 0x0628
    x"41",x"96",x"4E",x"B9",x"BA",x"02",x"C9",x"70", -- 0x0630
    x"F0",x"11",x"C9",x"A0",x"F0",x"07",x"8A",x"0A", -- 0x0638
    x"0A",x"0A",x"18",x"69",x"78",x"99",x"BA",x"02", -- 0x0640
    x"4C",x"31",x"A5",x"A4",x"01",x"B9",x"A2",x"02", -- 0x0648
    x"19",x"A3",x"02",x"29",x"02",x"F0",x"F1",x"4C", -- 0x0650
    x"5A",x"A5",x"A6",x"01",x"B5",x"51",x"DD",x"A2", -- 0x0658
    x"02",x"D0",x"06",x"A5",x"A2",x"29",x"01",x"F0", -- 0x0660
    x"10",x"38",x"FD",x"A2",x"02",x"B0",x"0A",x"A0", -- 0x0668
    x"02",x"84",x"61",x"A0",x"00",x"84",x"64",x"F0", -- 0x0670
    x"08",x"A0",x"00",x"84",x"61",x"A0",x"02",x"84", -- 0x0678
    x"64",x"B5",x"52",x"DD",x"A3",x"02",x"D0",x"06", -- 0x0680
    x"A5",x"A2",x"29",x"01",x"F0",x"10",x"38",x"FD", -- 0x0688
    x"A3",x"02",x"B0",x"0A",x"A0",x"03",x"84",x"62", -- 0x0690
    x"A0",x"01",x"84",x"63",x"D0",x"08",x"A0",x"01", -- 0x0698
    x"84",x"62",x"A0",x"03",x"84",x"63",x"A6",x"01", -- 0x06A0
    x"8A",x"0A",x"0A",x"0A",x"C5",x"A2",x"B0",x"2A", -- 0x06A8
    x"B5",x"51",x"38",x"FD",x"A2",x"02",x"B0",x"02", -- 0x06B0
    x"49",x"FF",x"85",x"69",x"B5",x"52",x"38",x"FD", -- 0x06B8
    x"A3",x"02",x"B0",x"02",x"49",x"FF",x"C5",x"69", -- 0x06C0
    x"90",x"10",x"A6",x"61",x"A4",x"62",x"86",x"62", -- 0x06C8
    x"84",x"61",x"A4",x"63",x"A6",x"64",x"84",x"64", -- 0x06D0
    x"86",x"63",x"A4",x"00",x"B9",x"BA",x"02",x"C9", -- 0x06D8
    x"A0",x"D0",x"08",x"A6",x"61",x"A4",x"63",x"86", -- 0x06E0
    x"63",x"84",x"61",x"60",x"A2",x"00",x"BD",x"F1", -- 0x06E8
    x"AB",x"9D",x"A2",x"02",x"E8",x"E0",x"0A",x"D0", -- 0x06F0
    x"F5",x"A0",x"00",x"BE",x"C4",x"AB",x"96",x"4B", -- 0x06F8
    x"C8",x"C0",x"10",x"D0",x"F6",x"60",x"E6",x"49", -- 0x0700
    x"A9",x"00",x"8D",x"A1",x"02",x"A9",x"0E",x"8D", -- 0x0708
    x"0F",x"90",x"A9",x"93",x"20",x"D2",x"FF",x"A2", -- 0x0710
    x"06",x"20",x"81",x"A7",x"A2",x"15",x"BD",x"00", -- 0x0718
    x"AC",x"9D",x"00",x"1E",x"BD",x"E3",x"AC",x"9D", -- 0x0720
    x"E3",x"1E",x"E8",x"D0",x"F1",x"86",x"4A",x"BD", -- 0x0728
    x"50",x"AE",x"9D",x"B2",x"02",x"A9",x"80",x"9D", -- 0x0730
    x"BA",x"02",x"A9",x"1C",x"9D",x"C2",x"02",x"E8", -- 0x0738
    x"E0",x"05",x"D0",x"EB",x"A4",x"45",x"20",x"AA", -- 0x0740
    x"AB",x"88",x"F0",x"0D",x"A9",x"19",x"99",x"E4", -- 0x0748
    x"1F",x"A9",x"07",x"99",x"E4",x"97",x"88",x"D0", -- 0x0750
    x"F3",x"A4",x"49",x"A2",x"00",x"C0",x"0C",x"90", -- 0x0758
    x"02",x"A0",x"0C",x"B9",x"55",x"AE",x"9D",x"F1", -- 0x0760
    x"1F",x"B9",x"62",x"AE",x"9D",x"F1",x"97",x"C0", -- 0x0768
    x"00",x"F0",x"0D",x"E8",x"86",x"FF",x"A5",x"49", -- 0x0770
    x"38",x"E5",x"FF",x"A8",x"E0",x"07",x"D0",x"DD", -- 0x0778
    x"60",x"A0",x"15",x"B9",x"00",x"AC",x"C9",x"29", -- 0x0780
    x"90",x"0A",x"C9",x"3F",x"B0",x"06",x"A9",x"01", -- 0x0788
    x"8A",x"99",x"00",x"96",x"B9",x"E3",x"AC",x"C9", -- 0x0790
    x"29",x"90",x"08",x"C9",x"3F",x"B0",x"04",x"8A", -- 0x0798
    x"99",x"E3",x"96",x"C8",x"D0",x"DD",x"60",x"A4", -- 0x07A0
    x"01",x"A5",x"40",x"29",x"01",x"F0",x"01",x"C8", -- 0x07A8
    x"B9",x"A2",x"02",x"29",x"07",x"F0",x"0E",x"A5", -- 0x07B0
    x"41",x"C5",x"40",x"F0",x"3C",x"45",x"40",x"C9", -- 0x07B8
    x"02",x"F0",x"36",x"38",x"60",x"20",x"76",x"A8", -- 0x07C0
    x"A5",x"F8",x"38",x"E9",x"04",x"85",x"F8",x"A6", -- 0x07C8
    x"41",x"E0",x"02",x"B0",x"0F",x"A5",x"F7",x"18", -- 0x07D0
    x"7D",x"E5",x"AB",x"90",x"02",x"E6",x"F8",x"85", -- 0x07D8
    x"F7",x"18",x"90",x"0C",x"A5",x"F7",x"38",x"FD", -- 0x07E0
    x"E3",x"AB",x"B0",x"02",x"C6",x"F8",x"85",x"F7", -- 0x07E8
    x"A0",x"00",x"B1",x"F7",x"C9",x"29",x"90",x"01", -- 0x07F0
    x"60",x"A5",x"41",x"0A",x"AA",x"A4",x"01",x"BD", -- 0x07F8
    x"DD",x"AB",x"18",x"79",x"A2",x"02",x"99",x"A2", -- 0x0800
    x"02",x"BD",x"DE",x"AB",x"18",x"79",x"A3",x"02", -- 0x0808
    x"99",x"A3",x"02",x"18",x"60",x"A9",x"00",x"85", -- 0x0810
    x"00",x"0A",x"85",x"01",x"0A",x"0A",x"85",x"02", -- 0x0818
    x"A6",x"00",x"AD",x"A1",x"02",x"3D",x"FB",x"AB", -- 0x0820
    x"F0",x"1A",x"AD",x"CC",x"02",x"3D",x"FB",x"AB", -- 0x0828
    x"F0",x"03",x"20",x"65",x"A8",x"20",x"76",x"A8", -- 0x0830
    x"20",x"E0",x"A8",x"20",x"3D",x"A9",x"20",x"E3", -- 0x0838
    x"A9",x"4C",x"4F",x"A8",x"AD",x"CC",x"02",x"3D", -- 0x0840
    x"FB",x"AB",x"F0",x"03",x"20",x"65",x"A8",x"E6", -- 0x0848
    x"00",x"A5",x"00",x"C9",x"05",x"D0",x"C2",x"A2", -- 0x0850
    x"00",x"BD",x"A1",x"02",x"9D",x"CC",x"02",x"E8", -- 0x0858
    x"E0",x"11",x"D0",x"F5",x"60",x"20",x"6F",x"A8", -- 0x0860
    x"20",x"E0",x"A8",x"20",x"18",x"A9",x"60",x"A5", -- 0x0868
    x"01",x"18",x"69",x"CC",x"D0",x"05",x"A5",x"01", -- 0x0870
    x"18",x"69",x"A1",x"AA",x"BD",x"01",x"02",x"C9", -- 0x0878
    x"A0",x"90",x"02",x"E9",x"A0",x"4A",x"4A",x"4A", -- 0x0880
    x"85",x"F7",x"85",x"FC",x"AD",x"88",x"02",x"85", -- 0x0888
    x"F8",x"A5",x"F4",x"29",x"FE",x"85",x"FD",x"BD", -- 0x0890
    x"02",x"02",x"C9",x"B8",x"90",x"02",x"E9",x"B8", -- 0x0898
    x"4A",x"4A",x"4A",x"A8",x"F0",x"12",x"A5",x"F7", -- 0x08A0
    x"18",x"69",x"15",x"90",x"04",x"E6",x"F8",x"E6", -- 0x08A8
    x"FD",x"85",x"F7",x"85",x"FC",x"88",x"D0",x"F0", -- 0x08B0
    x"A5",x"F8",x"85",x"FA",x"A5",x"FD",x"85",x"FF", -- 0x08B8
    x"BD",x"01",x"02",x"29",x"07",x"F0",x"10",x"A5", -- 0x08C0
    x"F7",x"18",x"69",x"01",x"90",x"04",x"E6",x"FA", -- 0x08C8
    x"E6",x"FF",x"85",x"F9",x"85",x"FE",x"60",x"A5", -- 0x08D0
    x"F7",x"18",x"69",x"15",x"90",x"F4",x"B0",x"EE", -- 0x08D8
    x"A0",x"00",x"B1",x"F7",x"48",x"A4",x"01",x"BD", -- 0x08E0
    x"01",x"02",x"29",x"07",x"D0",x"07",x"BD",x"02", -- 0x08E8
    x"02",x"29",x"07",x"F0",x"08",x"A0",x"00",x"B1", -- 0x08F0
    x"F9",x"48",x"A4",x"01",x"C8",x"98",x"AA",x"68", -- 0x08F8
    x"C5",x"01",x"90",x"0B",x"C9",x"0A",x"B0",x"07", -- 0x0900
    x"A8",x"B9",x"DD",x"02",x"18",x"90",x"F1",x"9D", -- 0x0908
    x"DD",x"02",x"CA",x"E4",x"01",x"F0",x"E8",x"60", -- 0x0910
    x"A6",x"01",x"BD",x"DD",x"02",x"A0",x"00",x"91", -- 0x0918
    x"F7",x"A9",x"01",x"91",x"FC",x"BD",x"CD",x"02", -- 0x0920
    x"29",x"07",x"D0",x"07",x"BD",x"CE",x"02",x"29", -- 0x0928
    x"07",x"F0",x"09",x"BD",x"DE",x"02",x"91",x"F9", -- 0x0930
    x"A9",x"01",x"91",x"FE",x"60",x"A6",x"00",x"BD", -- 0x0938
    x"BA",x"02",x"85",x"05",x"BD",x"C2",x"02",x"85", -- 0x0940
    x"06",x"A6",x"01",x"BD",x"A3",x"02",x"29",x"07", -- 0x0948
    x"85",x"03",x"AA",x"A0",x"00",x"98",x"99",x"5C", -- 0x0950
    x"03",x"C8",x"C0",x"10",x"D0",x"F8",x"A8",x"B1", -- 0x0958
    x"05",x"9D",x"5C",x"03",x"E8",x"C8",x"C0",x"08", -- 0x0960
    x"D0",x"F5",x"A6",x"01",x"BD",x"A2",x"02",x"29", -- 0x0968
    x"07",x"A8",x"F0",x"11",x"A2",x"00",x"18",x"7E", -- 0x0970
    x"5C",x"03",x"7E",x"64",x"03",x"E8",x"E0",x"08", -- 0x0978
    x"D0",x"F4",x"88",x"D0",x"EF",x"84",x"FB",x"A5", -- 0x0980
    x"01",x"18",x"65",x"FB",x"AA",x"A9",x"1C",x"85", -- 0x0988
    x"06",x"BD",x"DD",x"02",x"C9",x"80",x"90",x"04", -- 0x0990
    x"A0",x"80",x"84",x"06",x"29",x"1F",x"0A",x"0A", -- 0x0998
    x"0A",x"85",x"05",x"BD",x"DD",x"02",x"29",x"60", -- 0x09A0
    x"4A",x"4A",x"4A",x"4A",x"4A",x"18",x"65",x"06", -- 0x09A8
    x"85",x"06",x"A0",x"00",x"A5",x"FB",x"0A",x"0A", -- 0x09B0
    x"0A",x"AA",x"B1",x"05",x"9D",x"6C",x"03",x"E8", -- 0x09B8
    x"C8",x"C0",x"08",x"D0",x"F5",x"E6",x"FB",x"A5", -- 0x09C0
    x"FB",x"C9",x"02",x"D0",x"BA",x"A0",x"00",x"A5", -- 0x09C8
    x"02",x"0A",x"AA",x"B9",x"5C",x"03",x"19",x"6C", -- 0x09D0
    x"03",x"9D",x"00",x"1C",x"E8",x"C8",x"C0",x"10", -- 0x09D8
    x"D0",x"F1",x"60",x"A5",x"01",x"A0",x"00",x"91", -- 0x09E0
    x"F7",x"A6",x"00",x"BD",x"B2",x"02",x"91",x"FC", -- 0x09E8
    x"A6",x"01",x"BD",x"A2",x"02",x"29",x"07",x"D0", -- 0x09F0
    x"07",x"BD",x"A3",x"02",x"29",x"07",x"F0",x"08", -- 0x09F8
    x"B1",x"FC",x"91",x"FE",x"E8",x"8A",x"91",x"F9", -- 0x0A00
    x"60",x"D8",x"AD",x"DC",x"1E",x"C9",x"C5",x"D0", -- 0x0A08
    x"05",x"A9",x"09",x"8D",x"DC",x"96",x"A5",x"A2", -- 0x0A10
    x"29",x"07",x"D0",x"3B",x"A5",x"10",x"F0",x"37", -- 0x0A18
    x"C9",x"1F",x"B0",x"18",x"29",x"03",x"D0",x"14", -- 0x0A20
    x"A0",x"04",x"B9",x"BA",x"02",x"C9",x"A0",x"D0", -- 0x0A28
    x"08",x"B9",x"B2",x"02",x"49",x"07",x"99",x"B2", -- 0x0A30
    x"02",x"88",x"D0",x"EE",x"C6",x"10",x"D0",x"17", -- 0x0A38
    x"A0",x"04",x"B9",x"50",x"AE",x"99",x"B2",x"02", -- 0x0A40
    x"B9",x"BA",x"02",x"C9",x"70",x"F0",x"05",x"A9", -- 0x0A48
    x"98",x"99",x"BA",x"02",x"88",x"D0",x"EB",x"A5", -- 0x0A50
    x"46",x"C9",x"1E",x"D0",x"2E",x"A2",x"00",x"86", -- 0x0A58
    x"46",x"BD",x"F8",x"1C",x"5D",x"88",x"82",x"9D", -- 0x0A60
    x"F8",x"1C",x"E8",x"E0",x"08",x"D0",x"F2",x"A9", -- 0x0A68
    x"FE",x"4D",x"9F",x"1C",x"8D",x"9F",x"1C",x"8D", -- 0x0A70
    x"A7",x"1C",x"8D",x"8F",x"1C",x"8D",x"97",x"1C", -- 0x0A78
    x"A9",x"7F",x"4D",x"7F",x"1C",x"8D",x"7F",x"1C", -- 0x0A80
    x"8D",x"87",x"1C",x"E6",x"46",x"A5",x"45",x"D0", -- 0x0A88
    x"1E",x"A5",x"A2",x"F0",x"1A",x"A5",x"A1",x"29", -- 0x0A90
    x"03",x"D0",x"14",x"E6",x"48",x"A5",x"48",x"29", -- 0x0A98
    x"03",x"0A",x"A8",x"B9",x"CC",x"AB",x"8D",x"A2", -- 0x0AA0
    x"02",x"B9",x"CD",x"AB",x"8D",x"A3",x"02",x"A2", -- 0x0AA8
    x"00",x"BD",x"06",x"1A",x"DD",x"0F",x"1A",x"90", -- 0x0AB0
    x"14",x"D0",x"05",x"E8",x"E0",x"06",x"D0",x"F1", -- 0x0AB8
    x"A2",x"00",x"BD",x"06",x"1A",x"9D",x"0F",x"1A", -- 0x0AC0
    x"E8",x"E0",x"06",x"D0",x"F5",x"A2",x"14",x"BD", -- 0x0AC8
    x"00",x"1A",x"9D",x"00",x"1E",x"CA",x"10",x"F7", -- 0x0AD0
    x"A4",x"3F",x"F0",x"19",x"A6",x"3E",x"BD",x"00", -- 0x0AD8
    x"1A",x"C9",x"B9",x"F0",x"08",x"FE",x"00",x"1A", -- 0x0AE0
    x"88",x"D0",x"F1",x"F0",x"08",x"A9",x"B0",x"9D", -- 0x0AE8
    x"00",x"1A",x"CA",x"D0",x"E9",x"84",x"3F",x"A2", -- 0x0AF0
    x"00",x"A0",x"00",x"B5",x"4B",x"D0",x"2E",x"BD", -- 0x0AF8
    x"BB",x"02",x"C9",x"70",x"D0",x"0C",x"A9",x"50", -- 0x0B00
    x"99",x"53",x"00",x"A9",x"48",x"99",x"54",x"00", -- 0x0B08
    x"D0",x"1B",x"A5",x"4A",x"C9",x"A6",x"B0",x"09", -- 0x0B10
    x"BD",x"C4",x"AB",x"F0",x"04",x"C5",x"A2",x"D0", -- 0x0B18
    x"0C",x"AD",x"A2",x"02",x"99",x"53",x"00",x"AD", -- 0x0B20
    x"A3",x"02",x"99",x"54",x"00",x"C8",x"C8",x"E8", -- 0x0B28
    x"E0",x"04",x"D0",x"C7",x"A5",x"3D",x"F0",x"05", -- 0x0B30
    x"A9",x"91",x"8D",x"0C",x"90",x"A9",x"00",x"85", -- 0x0B38
    x"3D",x"AD",x"0C",x"90",x"F0",x"23",x"AD",x"0C", -- 0x0B40
    x"90",x"29",x"01",x"F0",x"13",x"AD",x"0C",x"90", -- 0x0B48
    x"18",x"69",x"10",x"C9",x"F1",x"90",x"03",x"38", -- 0x0B50
    x"E9",x"01",x"8D",x"0C",x"90",x"18",x"90",x"09", -- 0x0B58
    x"AD",x"0C",x"90",x"38",x"E9",x"10",x"8D",x"0C", -- 0x0B60
    x"90",x"A6",x"3C",x"F0",x"0E",x"A5",x"A2",x"29", -- 0x0B68
    x"01",x"D0",x"08",x"BD",x"E7",x"AB",x"8D",x"0B", -- 0x0B70
    x"90",x"C6",x"3C",x"A5",x"47",x"D0",x"17",x"AD", -- 0x0B78
    x"07",x"1A",x"C9",x"B1",x"D0",x"10",x"85",x"47", -- 0x0B80
    x"A6",x"45",x"A9",x"19",x"9D",x"E4",x"1F",x"A9", -- 0x0B88
    x"07",x"9D",x"E4",x"97",x"E6",x"45",x"4C",x"BF", -- 0x0B90
    x"EA",x"48",x"8A",x"48",x"20",x"15",x"A8",x"68", -- 0x0B98
    x"AA",x"68",x"18",x"65",x"A2",x"C5",x"A2",x"D0", -- 0x0BA0
    x"FC",x"60",x"A2",x"08",x"BD",x"D4",x"AB",x"C0", -- 0x0BA8
    x"00",x"F0",x"02",x"A9",x"20",x"9D",x"17",x"1F", -- 0x0BB0
    x"9D",x"17",x"1B",x"A9",x"02",x"9D",x"17",x"97", -- 0x0BB8
    x"CA",x"10",x"E9",x"60",x"00",x"33",x"76",x"F9", -- 0x0BC0
    x"00",x"03",x"02",x"00",x"A0",x"28",x"00",x"28", -- 0x0BC8
    x"A0",x"88",x"00",x"88",x"87",x"81",x"8D",x"85", -- 0x0BD0
    x"A0",x"8F",x"96",x"85",x"92",x"01",x"00",x"00", -- 0x0BD8
    x"01",x"FF",x"00",x"00",x"FF",x"01",x"15",x"00", -- 0x0BE0
    x"00",x"C0",x"B8",x"B0",x"A8",x"B0",x"B8",x"C0", -- 0x0BE8
    x"C8",x"50",x"88",x"50",x"48",x"50",x"58",x"60", -- 0x0BF0
    x"58",x"40",x"58",x"01",x"02",x"04",x"08",x"10", -- 0x0BF8
    x"93",x"83",x"8F",x"92",x"85",x"BA",x"B0",x"B0", -- 0x0C00
    x"B0",x"B0",x"B0",x"B0",x"A0",x"A0",x"A0",x"B0", -- 0x0C08
    x"B2",x"B0",x"B0",x"B0",x"B0",x"37",x"3A",x"3A", -- 0x0C10
    x"3A",x"3A",x"3A",x"3A",x"3A",x"3A",x"3A",x"3D", -- 0x0C18
    x"3A",x"3A",x"3A",x"3A",x"3A",x"3A",x"3A",x"3A", -- 0x0C20
    x"3A",x"38",x"39",x"1E",x"1E",x"1E",x"1E",x"1E", -- 0x0C28
    x"1E",x"1E",x"1E",x"1E",x"39",x"1E",x"1E",x"1E", -- 0x0C30
    x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"39",x"39", -- 0x0C38
    x"1E",x"2F",x"30",x"1E",x"2F",x"2B",x"2B",x"30", -- 0x0C40
    x"1E",x"39",x"1E",x"2F",x"2B",x"2B",x"30",x"1E", -- 0x0C48
    x"2F",x"30",x"1E",x"39",x"39",x"1F",x"2D",x"2E", -- 0x0C50
    x"1E",x"2D",x"2C",x"2C",x"2E",x"1E",x"32",x"1E", -- 0x0C58
    x"2D",x"2C",x"2C",x"2E",x"1E",x"2D",x"2E",x"1F", -- 0x0C60
    x"39",x"39",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E", -- 0x0C68
    x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E", -- 0x0C70
    x"1E",x"1E",x"1E",x"1E",x"1E",x"39",x"39",x"1E", -- 0x0C78
    x"33",x"34",x"1E",x"31",x"1E",x"33",x"3A",x"3A", -- 0x0C80
    x"3D",x"3A",x"3A",x"34",x"1E",x"31",x"1E",x"33", -- 0x0C88
    x"34",x"1E",x"39",x"39",x"1E",x"1E",x"1E",x"1E", -- 0x0C90
    x"39",x"1E",x"1E",x"1E",x"1E",x"39",x"1E",x"1E", -- 0x0C98
    x"1E",x"1E",x"39",x"1E",x"1E",x"1E",x"1E",x"39", -- 0x0CA0
    x"35",x"3A",x"3A",x"38",x"1E",x"3B",x"3A",x"3A", -- 0x0CA8
    x"34",x"20",x"32",x"20",x"33",x"3A",x"3A",x"3C", -- 0x0CB0
    x"1E",x"37",x"3A",x"3A",x"36",x"20",x"20",x"20", -- 0x0CB8
    x"39",x"1E",x"39",x"20",x"20",x"20",x"20",x"20", -- 0x0CC0
    x"20",x"20",x"20",x"20",x"39",x"1E",x"39",x"20", -- 0x0CC8
    x"20",x"20",x"3A",x"3A",x"3A",x"36",x"1E",x"32", -- 0x0CD0
    x"20",x"37",x"3A",x"29",x"C5",x"2A",x"3A",x"38", -- 0x0CD8
    x"20",x"32",x"1E",x"35",x"3A",x"3A",x"3A",x"20", -- 0x0CE0
    x"20",x"20",x"20",x"1E",x"20",x"20",x"39",x"20", -- 0x0CE8
    x"20",x"20",x"20",x"20",x"39",x"20",x"20",x"1E", -- 0x0CF0
    x"20",x"20",x"20",x"20",x"3A",x"3A",x"3A",x"38", -- 0x0CF8
    x"1E",x"31",x"20",x"35",x"3A",x"3A",x"3A",x"3A", -- 0x0D00
    x"3A",x"36",x"20",x"31",x"1E",x"37",x"3A",x"3A", -- 0x0D08
    x"3A",x"20",x"20",x"20",x"39",x"1E",x"39",x"20", -- 0x0D10
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x0D18
    x"39",x"1E",x"39",x"20",x"20",x"20",x"37",x"3A", -- 0x0D20
    x"3A",x"36",x"1E",x"32",x"20",x"33",x"3A",x"3A", -- 0x0D28
    x"3D",x"3A",x"3A",x"34",x"20",x"32",x"1E",x"35", -- 0x0D30
    x"3A",x"3A",x"38",x"39",x"1E",x"1E",x"1E",x"1E", -- 0x0D38
    x"1E",x"1E",x"1E",x"1E",x"1E",x"39",x"1E",x"1E", -- 0x0D40
    x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"39", -- 0x0D48
    x"39",x"1E",x"33",x"38",x"1E",x"33",x"3A",x"3A", -- 0x0D50
    x"34",x"1E",x"32",x"1E",x"33",x"3A",x"3A",x"34", -- 0x0D58
    x"1E",x"37",x"34",x"1E",x"39",x"39",x"1F",x"1E", -- 0x0D60
    x"39",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"20", -- 0x0D68
    x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"39",x"1E", -- 0x0D70
    x"1F",x"39",x"3B",x"34",x"1E",x"32",x"1E",x"31", -- 0x0D78
    x"1E",x"33",x"3A",x"3A",x"3D",x"3A",x"3A",x"34", -- 0x0D80
    x"1E",x"31",x"1E",x"32",x"1E",x"33",x"3C",x"39", -- 0x0D88
    x"1E",x"1E",x"1E",x"1E",x"39",x"1E",x"1E",x"1E", -- 0x0D90
    x"1E",x"39",x"1E",x"1E",x"1E",x"1E",x"39",x"1E", -- 0x0D98
    x"1E",x"1E",x"1E",x"39",x"39",x"1E",x"33",x"3A", -- 0x0DA0
    x"3A",x"3E",x"3A",x"3A",x"34",x"1E",x"32",x"1E", -- 0x0DA8
    x"33",x"3A",x"3A",x"3E",x"3A",x"3A",x"34",x"1E", -- 0x0DB0
    x"39",x"39",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E", -- 0x0DB8
    x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E", -- 0x0DC0
    x"1E",x"1E",x"1E",x"1E",x"1E",x"39",x"35",x"3A", -- 0x0DC8
    x"3A",x"3A",x"3A",x"3A",x"3A",x"3A",x"3A",x"3A", -- 0x0DD0
    x"3A",x"3A",x"3A",x"3A",x"3A",x"3A",x"3A",x"3A", -- 0x0DD8
    x"3A",x"3A",x"36",x"3F",x"B2",x"B0",x"B0",x"B8", -- 0x0DE0
    x"A0",x"92",x"88",x"95",x"92",x"93",x"94",x"A0", -- 0x0DE8
    x"A0",x"00",x"01",x"93",x"94",x"81",x"92",x"94", -- 0x0DF0
    x"01",x"03",x"05",x"07",x"0A",x"14",x"1E",x"32", -- 0x0DF8
    x"FF",x"EA",x"EF",x"EF",x"EB",x"EF",x"EF",x"FF", -- 0x0E00
    x"FC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"FC", -- 0x0E08
    x"38",x"7C",x"FE",x"92",x"FE",x"FE",x"FE",x"AA", -- 0x0E10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E18
    x"38",x"7C",x"FE",x"92",x"FE",x"FE",x"FE",x"AA", -- 0x0E20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E28
    x"38",x"7C",x"FE",x"92",x"FE",x"FE",x"FE",x"AA", -- 0x0E30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E38
    x"38",x"7C",x"FE",x"92",x"FE",x"FE",x"FE",x"AA", -- 0x0E40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E48
    x"07",x"02",x"05",x"03",x"07",x"21",x"22",x"23", -- 0x0E50
    x"23",x"24",x"24",x"25",x"25",x"26",x"26",x"27", -- 0x0E58
    x"27",x"28",x"02",x"02",x"07",x"07",x"02",x"02", -- 0x0E60
    x"05",x"05",x"04",x"04",x"07",x"07",x"03",x"00", -- 0x0E68
    x"00",x"38",x"7C",x"54",x"7C",x"7C",x"54",x"00", -- 0x0E70
    x"1C",x"3E",x"7F",x"64",x"7F",x"7F",x"7F",x"55", -- 0x0E78
    x"1C",x"3E",x"7F",x"7F",x"49",x"7F",x"7F",x"55", -- 0x0E80
    x"38",x"7C",x"FE",x"26",x"FE",x"FE",x"FE",x"AA", -- 0x0E88
    x"38",x"7C",x"FE",x"FE",x"FE",x"FE",x"FE",x"AA", -- 0x0E90
    x"38",x"7C",x"FE",x"92",x"FE",x"82",x"FE",x"AA", -- 0x0E98
    x"38",x"7C",x"FE",x"92",x"FE",x"82",x"FE",x"54", -- 0x0EA0
    x"3C",x"7E",x"BD",x"FF",x"BD",x"C3",x"7E",x"3C", -- 0x0EA8
    x"3C",x"7E",x"FF",x"FF",x"FF",x"FF",x"7E",x"3C", -- 0x0EB0
    x"3E",x"7C",x"F8",x"F0",x"F0",x"F8",x"7C",x"3E", -- 0x0EB8
    x"3C",x"7E",x"FF",x"FF",x"E7",x"C3",x"81",x"00", -- 0x0EC0
    x"7C",x"3E",x"1F",x"0F",x"0F",x"1F",x"3E",x"7C", -- 0x0EC8
    x"00",x"81",x"C3",x"E7",x"FF",x"FF",x"7E",x"3C", -- 0x0ED0
    x"00",x"10",x"10",x"6C",x"10",x"10",x"00",x"00", -- 0x0ED8
    x"10",x"44",x"28",x"C6",x"28",x"44",x"10",x"00", -- 0x0EE0
    x"92",x"44",x"00",x"82",x"00",x"44",x"92",x"00", -- 0x0EE8
    x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00", -- 0x0EF0
    x"00",x"3C",x"7E",x"7E",x"7E",x"7E",x"3C",x"00", -- 0x0EF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F00
    x"04",x"08",x"18",x"24",x"62",x"F7",x"F2",x"60", -- 0x0F08
    x"10",x"7C",x"FE",x"AA",x"D6",x"AA",x"54",x"28", -- 0x0F10
    x"20",x"10",x"7C",x"FE",x"FE",x"FE",x"7C",x"38", -- 0x0F18
    x"08",x"10",x"7C",x"FE",x"FE",x"FE",x"7C",x"28", -- 0x0F20
    x"08",x"10",x"38",x"38",x"7C",x"FE",x"FE",x"6C", -- 0x0F28
    x"10",x"30",x"92",x"FE",x"7C",x"38",x"10",x"28", -- 0x0F30
    x"10",x"38",x"7C",x"7C",x"7C",x"7C",x"FE",x"10", -- 0x0F38
    x"18",x"24",x"18",x"08",x"08",x"18",x"08",x"18", -- 0x0F40
    x"00",x"FF",x"01",x"01",x"01",x"01",x"FE",x"00", -- 0x0F48
    x"00",x"FF",x"80",x"80",x"80",x"80",x"7F",x"00", -- 0x0F50
    x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F58
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00", -- 0x0F60
    x"40",x"40",x"40",x"40",x"40",x"20",x"1F",x"00", -- 0x0F68
    x"02",x"02",x"02",x"02",x"02",x"04",x"F8",x"00", -- 0x0F70
    x"00",x"1F",x"20",x"40",x"40",x"40",x"40",x"40", -- 0x0F78
    x"00",x"F8",x"04",x"02",x"02",x"02",x"02",x"02", -- 0x0F80
    x"00",x"18",x"24",x"42",x"42",x"42",x"42",x"42", -- 0x0F88
    x"42",x"42",x"42",x"42",x"42",x"24",x"18",x"00", -- 0x0F90
    x"00",x"1F",x"20",x"40",x"40",x"20",x"1F",x"00", -- 0x0F98
    x"00",x"F8",x"04",x"02",x"02",x"04",x"F8",x"00", -- 0x0FA0
    x"42",x"41",x"40",x"40",x"40",x"20",x"1F",x"00", -- 0x0FA8
    x"42",x"82",x"02",x"02",x"02",x"04",x"F8",x"00", -- 0x0FB0
    x"00",x"1F",x"20",x"40",x"40",x"40",x"41",x"42", -- 0x0FB8
    x"00",x"F8",x"04",x"02",x"02",x"02",x"82",x"42", -- 0x0FC0
    x"42",x"42",x"42",x"42",x"42",x"42",x"42",x"42", -- 0x0FC8
    x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00", -- 0x0FD0
    x"42",x"41",x"40",x"40",x"40",x"40",x"41",x"42", -- 0x0FD8
    x"42",x"82",x"02",x"02",x"02",x"02",x"82",x"42", -- 0x0FE0
    x"00",x"FF",x"00",x"00",x"00",x"00",x"81",x"42", -- 0x0FE8
    x"42",x"81",x"00",x"00",x"00",x"00",x"FF",x"00", -- 0x0FF0
    x"3C",x"42",x"99",x"A1",x"A1",x"99",x"42",x"3C", -- 0x0FF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1000
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1008
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1010
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1018
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1020
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1028
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1030
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1038
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1040
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1048
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1050
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1058
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1060
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1068
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1070
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1078
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1080
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1088
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1090
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1098
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1100
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1108
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1110
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1118
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1120
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1128
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1130
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1138
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1140
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1148
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1150
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1158
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1160
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1168
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1170
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1178
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1180
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1188
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1190
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1198
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1200
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1208
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1210
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1218
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1220
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1228
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1230
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1238
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1240
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1248
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1250
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1258
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1260
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1268
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1270
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1278
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1280
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1288
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1290
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1298
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1300
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1308
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1310
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1318
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1320
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1328
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1330
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1338
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1340
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1348
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1350
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1358
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1360
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1368
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1370
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1378
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1380
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1388
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1390
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1398
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1400
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1408
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1410
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1418
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1420
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1428
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1430
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1438
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1440
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1448
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1450
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1458
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1460
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1468
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1470
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1478
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1480
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1488
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1490
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1498
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1500
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1508
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1510
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1518
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1520
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1528
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1530
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1538
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1540
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1548
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1550
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1558
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1560
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1568
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1570
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1578
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1580
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1588
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1590
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1598
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1600
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1608
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1610
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1618
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1620
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1628
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1630
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1638
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1640
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1648
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1650
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1658
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1660
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1668
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1670
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1678
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1680
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1688
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1690
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1698
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1700
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1708
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1710
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1718
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1720
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1728
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1730
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1738
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1740
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1748
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1750
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1758
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1760
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1768
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1770
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1778
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1780
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1788
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1790
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1798
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1800
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1808
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1810
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1818
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1820
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1828
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1830
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1838
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1840
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1848
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1850
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1858
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1860
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1868
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1870
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1878
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1880
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1888
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1890
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1898
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1900
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1908
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1910
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1918
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1920
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1928
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1930
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1938
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1940
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1948
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1950
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1958
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1960
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1968
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1970
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1978
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1980
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1988
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1990
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1998
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x1FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
