-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity cart_rom is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of cart_rom is


  type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"D5",x"A8",x"09",x"A0",x"41",x"30",x"C3",x"C2", -- 0x0000
    x"CD",x"68",x"A8",x"68",x"AA",x"68",x"40",x"00", -- 0x0008
    x"BB",x"A2",x"AE",x"A7",x"C4",x"A7",x"8C",x"A1", -- 0x0010
    x"D5",x"A8",x"96",x"A8",x"16",x"A8",x"E1",x"A7", -- 0x0018
    x"0C",x"A5",x"A8",x"A8",x"B8",x"A5",x"80",x"A6", -- 0x0020
    x"22",x"A7",x"34",x"A2",x"82",x"A3",x"8F",x"A3", -- 0x0028
    x"A3",x"A3",x"AD",x"A3",x"4A",x"A0",x"17",x"A4", -- 0x0030
    x"52",x"A4",x"81",x"A4",x"91",x"A4",x"03",x"A8", -- 0x0038
    x"DB",x"A4",x"E0",x"A4",x"98",x"A1",x"A3",x"A5", -- 0x0040
    x"E5",x"A4",x"85",x"7F",x"86",x"76",x"84",x"77", -- 0x0048
    x"A2",x"2F",x"A9",x"00",x"95",x"BF",x"CA",x"10", -- 0x0050
    x"FB",x"A5",x"76",x"AA",x"4A",x"4A",x"4A",x"48", -- 0x0058
    x"8A",x"29",x"07",x"48",x"A9",x"00",x"85",x"71", -- 0x0060
    x"A5",x"7F",x"0A",x"0A",x"0A",x"0A",x"26",x"71", -- 0x0068
    x"69",x"D1",x"85",x"70",x"A5",x"71",x"69",x"AA", -- 0x0070
    x"85",x"71",x"A0",x"0F",x"B1",x"70",x"99",x"BF", -- 0x0078
    x"00",x"88",x"10",x"F8",x"68",x"F0",x"44",x"AA", -- 0x0080
    x"46",x"BF",x"66",x"D7",x"46",x"C0",x"66",x"D8", -- 0x0088
    x"46",x"C1",x"66",x"D9",x"46",x"C2",x"66",x"DA", -- 0x0090
    x"46",x"C3",x"66",x"DB",x"46",x"C4",x"66",x"DC", -- 0x0098
    x"46",x"C5",x"66",x"DD",x"46",x"C6",x"66",x"DE", -- 0x00A0
    x"46",x"C7",x"66",x"DF",x"46",x"C8",x"66",x"E0", -- 0x00A8
    x"46",x"C9",x"66",x"E1",x"46",x"CA",x"66",x"E2", -- 0x00B0
    x"46",x"CB",x"66",x"E3",x"46",x"CC",x"66",x"E4", -- 0x00B8
    x"46",x"CD",x"66",x"E5",x"46",x"CE",x"66",x"E6", -- 0x00C0
    x"CA",x"D0",x"BD",x"A5",x"77",x"A8",x"4A",x"4A", -- 0x00C8
    x"4A",x"48",x"98",x"29",x"07",x"F0",x"1F",x"18", -- 0x00D0
    x"69",x"0F",x"A8",x"A2",x"0F",x"B5",x"BF",x"99", -- 0x00D8
    x"BF",x"00",x"B5",x"D7",x"99",x"D7",x"00",x"88", -- 0x00E0
    x"CA",x"10",x"F2",x"A9",x"00",x"99",x"BF",x"00", -- 0x00E8
    x"99",x"D7",x"00",x"88",x"10",x"F7",x"A6",x"92", -- 0x00F0
    x"86",x"73",x"A4",x"93",x"84",x"74",x"20",x"96", -- 0x00F8
    x"A7",x"A9",x"45",x"85",x"72",x"A2",x"05",x"BC", -- 0x0100
    x"94",x"A9",x"B1",x"6E",x"C5",x"72",x"D0",x"06", -- 0x0108
    x"B5",x"9B",x"F0",x"02",x"91",x"6E",x"C6",x"72", -- 0x0110
    x"CA",x"10",x"EC",x"68",x"85",x"74",x"85",x"93", -- 0x0118
    x"68",x"85",x"73",x"85",x"92",x"20",x"96",x"A7", -- 0x0120
    x"A9",x"05",x"85",x"75",x"A6",x"75",x"A9",x"00", -- 0x0128
    x"95",x"8C",x"85",x"71",x"BC",x"94",x"A9",x"B1", -- 0x0130
    x"6E",x"95",x"9B",x"0A",x"26",x"71",x"0A",x"26", -- 0x0138
    x"71",x"0A",x"26",x"71",x"69",x"00",x"85",x"70", -- 0x0140
    x"A5",x"71",x"69",x"10",x"85",x"71",x"8A",x"0A", -- 0x0148
    x"0A",x"0A",x"AA",x"86",x"72",x"A0",x"00",x"B1", -- 0x0150
    x"70",x"35",x"BF",x"D0",x"08",x"E8",x"C8",x"C0", -- 0x0158
    x"08",x"D0",x"F4",x"F0",x"06",x"A6",x"75",x"B5", -- 0x0160
    x"9B",x"95",x"8C",x"A6",x"72",x"A0",x"00",x"B1", -- 0x0168
    x"70",x"15",x"BF",x"9D",x"00",x"12",x"E8",x"C8", -- 0x0170
    x"C0",x"08",x"D0",x"F3",x"A6",x"75",x"BC",x"94", -- 0x0178
    x"A9",x"8A",x"18",x"69",x"40",x"91",x"6E",x"C6", -- 0x0180
    x"75",x"10",x"A1",x"60",x"A8",x"20",x"A4",x"AE", -- 0x0188
    x"49",x"FF",x"4A",x"18",x"69",x"08",x"85",x"68", -- 0x0190
    x"86",x"95",x"C9",x"08",x"B0",x"04",x"A9",x"08", -- 0x0198
    x"D0",x"06",x"C9",x"88",x"90",x"02",x"A9",x"87", -- 0x01A0
    x"48",x"4A",x"4A",x"4A",x"85",x"69",x"68",x"29", -- 0x01A8
    x"07",x"85",x"72",x"A4",x"95",x"D0",x"03",x"A2", -- 0x01B0
    x"00",x"2C",x"A2",x"38",x"A0",x"00",x"BD",x"61", -- 0x01B8
    x"AA",x"99",x"BF",x"00",x"E8",x"C8",x"C0",x"38", -- 0x01C0
    x"D0",x"F4",x"C6",x"72",x"30",x"15",x"A2",x"07", -- 0x01C8
    x"56",x"BF",x"76",x"C7",x"56",x"CF",x"76",x"D7", -- 0x01D0
    x"76",x"DF",x"76",x"E7",x"76",x"EF",x"CA",x"10", -- 0x01D8
    x"EF",x"30",x"E7",x"A6",x"94",x"D0",x"01",x"E8", -- 0x01E0
    x"A9",x"20",x"9D",x"10",x"1A",x"9D",x"11",x"1A", -- 0x01E8
    x"9D",x"13",x"1A",x"9D",x"14",x"1A",x"A0",x"05", -- 0x01F0
    x"9D",x"26",x"1A",x"E8",x"88",x"D0",x"F9",x"A2", -- 0x01F8
    x"37",x"B5",x"BF",x"9D",x"A0",x"12",x"CA",x"10", -- 0x0200
    x"F8",x"A6",x"69",x"86",x"94",x"A9",x"54",x"18", -- 0x0208
    x"A4",x"95",x"D0",x"0A",x"9D",x"10",x"1A",x"69", -- 0x0210
    x"01",x"9D",x"11",x"1A",x"90",x"08",x"9D",x"13", -- 0x0218
    x"1A",x"69",x"01",x"9D",x"14",x"1A",x"69",x"01", -- 0x0220
    x"A0",x"05",x"9D",x"26",x"1A",x"E8",x"69",x"01", -- 0x0228
    x"88",x"D0",x"F7",x"60",x"A9",x"03",x"85",x"74", -- 0x0230
    x"A9",x"00",x"85",x"73",x"A2",x"00",x"86",x"7D", -- 0x0238
    x"A5",x"88",x"F0",x"04",x"C6",x"88",x"D0",x"72", -- 0x0240
    x"A9",x"05",x"85",x"88",x"20",x"96",x"A7",x"A9", -- 0x0248
    x"0A",x"85",x"72",x"A4",x"7D",x"B9",x"98",x"00", -- 0x0250
    x"C0",x"01",x"F0",x"0B",x"18",x"69",x"01",x"C9", -- 0x0258
    x"A8",x"D0",x"0D",x"A9",x"08",x"D0",x"09",x"38", -- 0x0260
    x"E9",x"01",x"C9",x"07",x"D0",x"02",x"A9",x"A7", -- 0x0268
    x"99",x"98",x"00",x"48",x"29",x"07",x"0A",x"09", -- 0x0270
    x"60",x"85",x"7E",x"68",x"4A",x"4A",x"4A",x"A8", -- 0x0278
    x"A6",x"7D",x"BD",x"9A",x"A9",x"AA",x"B5",x"A1", -- 0x0280
    x"D0",x"04",x"A9",x"20",x"D0",x"02",x"A5",x"7E", -- 0x0288
    x"91",x"6E",x"C8",x"C0",x"15",x"D0",x"02",x"A0", -- 0x0290
    x"01",x"C9",x"20",x"F0",x"03",x"18",x"69",x"01", -- 0x0298
    x"91",x"6E",x"C8",x"C0",x"15",x"D0",x"02",x"A0", -- 0x02A0
    x"01",x"E8",x"C6",x"72",x"D0",x"D8",x"E6",x"74", -- 0x02A8
    x"E6",x"74",x"E6",x"7D",x"A5",x"7D",x"C9",x"03", -- 0x02B0
    x"D0",x"92",x"60",x"85",x"72",x"F0",x"04",x"A9", -- 0x02B8
    x"08",x"D0",x"15",x"A5",x"80",x"F0",x"05",x"C6", -- 0x02C0
    x"80",x"4C",x"DA",x"A2",x"A9",x"0A",x"85",x"80", -- 0x02C8
    x"E6",x"81",x"A5",x"81",x"29",x"03",x"85",x"81", -- 0x02D0
    x"85",x"7F",x"20",x"4C",x"A0",x"A9",x"00",x"85", -- 0x02D8
    x"68",x"85",x"69",x"85",x"6A",x"A9",x"05",x"85", -- 0x02E0
    x"75",x"A6",x"75",x"B5",x"8C",x"C9",x"5B",x"F0", -- 0x02E8
    x"04",x"C9",x"54",x"B0",x"08",x"C5",x"68",x"90", -- 0x02F0
    x"4F",x"85",x"68",x"B0",x"4B",x"C9",x"60",x"90", -- 0x02F8
    x"47",x"A9",x"60",x"85",x"68",x"8A",x"C9",x"03", -- 0x0300
    x"08",x"90",x"02",x"E9",x"03",x"18",x"65",x"74", -- 0x0308
    x"38",x"E9",x"03",x"4A",x"AA",x"B5",x"98",x"4A", -- 0x0310
    x"4A",x"4A",x"85",x"72",x"A5",x"73",x"28",x"90", -- 0x0318
    x"03",x"18",x"69",x"01",x"38",x"E5",x"72",x"B0", -- 0x0320
    x"02",x"69",x"14",x"4A",x"18",x"7D",x"9A",x"A9", -- 0x0328
    x"A8",x"B9",x"A1",x"00",x"F0",x"12",x"BD",x"9D", -- 0x0330
    x"A9",x"18",x"65",x"69",x"85",x"69",x"A9",x"00", -- 0x0338
    x"99",x"A1",x"00",x"E6",x"6A",x"20",x"8F",x"A3", -- 0x0340
    x"C6",x"75",x"10",x"9D",x"A0",x"02",x"BE",x"9A", -- 0x0348
    x"A9",x"A9",x"0A",x"85",x"75",x"A9",x"00",x"15", -- 0x0350
    x"A1",x"E8",x"C6",x"75",x"D0",x"F9",x"49",x"FF", -- 0x0358
    x"99",x"6B",x"00",x"F0",x"03",x"20",x"6C",x"A3", -- 0x0360
    x"88",x"10",x"E3",x"60",x"8A",x"48",x"98",x"48", -- 0x0368
    x"BE",x"9A",x"A9",x"A0",x"0A",x"A9",x"FF",x"95", -- 0x0370
    x"A1",x"E8",x"88",x"D0",x"FA",x"68",x"A8",x"68", -- 0x0378
    x"AA",x"60",x"A5",x"97",x"F0",x"08",x"A9",x"10", -- 0x0380
    x"85",x"82",x"A9",x"01",x"85",x"83",x"60",x"A5", -- 0x0388
    x"97",x"F0",x"0F",x"A9",x"10",x"85",x"84",x"A9", -- 0x0390
    x"01",x"85",x"85",x"A9",x"00",x"85",x"82",x"8D", -- 0x0398
    x"0A",x"90",x"60",x"A9",x"10",x"85",x"86",x"A9", -- 0x03A0
    x"01",x"85",x"87",x"D0",x"EE",x"A5",x"82",x"F0", -- 0x03A8
    x"19",x"C6",x"83",x"D0",x"15",x"A9",x"02",x"85", -- 0x03B0
    x"83",x"C6",x"82",x"A5",x"82",x"48",x"8D",x"0E", -- 0x03B8
    x"90",x"18",x"69",x"80",x"8D",x"0A",x"90",x"68", -- 0x03C0
    x"F0",x"D1",x"A5",x"84",x"F0",x"1B",x"C6",x"85", -- 0x03C8
    x"D0",x"17",x"A9",x"01",x"85",x"85",x"A9",x"EE", -- 0x03D0
    x"8D",x"0D",x"90",x"C6",x"84",x"C6",x"84",x"A5", -- 0x03D8
    x"84",x"8D",x"0E",x"90",x"D0",x"03",x"8D",x"0D", -- 0x03E0
    x"90",x"A5",x"86",x"F0",x"29",x"C6",x"87",x"D0", -- 0x03E8
    x"25",x"A9",x"03",x"85",x"87",x"C6",x"86",x"A5", -- 0x03F0
    x"97",x"F0",x"1B",x"A5",x"86",x"85",x"72",x"A9", -- 0x03F8
    x"0F",x"38",x"E5",x"72",x"8D",x"0E",x"90",x"A5", -- 0x0400
    x"72",x"18",x"69",x"BB",x"8D",x"0C",x"90",x"A5", -- 0x0408
    x"86",x"D0",x"03",x"8D",x"0C",x"90",x"60",x"AA", -- 0x0410
    x"BD",x"5E",x"AA",x"AA",x"A9",x"00",x"8D",x"0A", -- 0x0418
    x"90",x"8D",x"0B",x"90",x"8D",x"0C",x"90",x"8D", -- 0x0420
    x"0D",x"90",x"A9",x"08",x"8D",x"0E",x"90",x"BD", -- 0x0428
    x"05",x"AA",x"F0",x"1A",x"8D",x"0C",x"90",x"BD", -- 0x0430
    x"06",x"AA",x"E8",x"E8",x"A8",x"C0",x"01",x"D0", -- 0x0438
    x"05",x"A9",x"00",x"8D",x"0C",x"90",x"20",x"96", -- 0x0440
    x"A8",x"88",x"D0",x"F1",x"F0",x"E1",x"8D",x"0E", -- 0x0448
    x"90",x"60",x"0A",x"0A",x"AA",x"A0",x"00",x"BD", -- 0x0450
    x"E6",x"A9",x"99",x"56",x"19",x"E8",x"C8",x"C0", -- 0x0458
    x"04",x"D0",x"F4",x"A2",x"04",x"BD",x"DC",x"A9", -- 0x0460
    x"9D",x"50",x"19",x"CA",x"10",x"F7",x"A9",x"01", -- 0x0468
    x"20",x"17",x"A4",x"A2",x"09",x"A9",x"20",x"9D", -- 0x0470
    x"24",x"19",x"9D",x"50",x"19",x"CA",x"10",x"F7", -- 0x0478
    x"60",x"A2",x"09",x"BD",x"DC",x"A9",x"9D",x"24", -- 0x0480
    x"19",x"CA",x"10",x"F7",x"A9",x"00",x"4C",x"17", -- 0x0488
    x"A4",x"48",x"8A",x"48",x"98",x"48",x"20",x"A3", -- 0x0490
    x"A3",x"20",x"34",x"A2",x"68",x"48",x"AA",x"A0", -- 0x0498
    x"B8",x"20",x"4C",x"A0",x"20",x"AD",x"A3",x"20", -- 0x04A0
    x"96",x"A8",x"A5",x"87",x"C9",x"03",x"D0",x"E9", -- 0x04A8
    x"A5",x"86",x"F0",x"0C",x"C9",x"0A",x"F0",x"04", -- 0x04B0
    x"C9",x"05",x"D0",x"DD",x"E6",x"7F",x"D0",x"D9", -- 0x04B8
    x"68",x"68",x"AA",x"68",x"A4",x"97",x"F0",x"12", -- 0x04C0
    x"20",x"03",x"A8",x"A9",x"02",x"20",x"17",x"A4", -- 0x04C8
    x"A2",x"0F",x"A9",x"20",x"9D",x"4D",x"19",x"CA", -- 0x04D0
    x"10",x"FA",x"60",x"A9",x"FF",x"85",x"97",x"60", -- 0x04D8
    x"A9",x"00",x"85",x"97",x"60",x"A5",x"8A",x"F0", -- 0x04E0
    x"03",x"C6",x"8A",x"60",x"A9",x"32",x"85",x"8A", -- 0x04E8
    x"A2",x"08",x"AD",x"24",x"19",x"C9",x"20",x"F0", -- 0x04F0
    x"09",x"A9",x"20",x"9D",x"24",x"19",x"CA",x"10", -- 0x04F8
    x"FA",x"60",x"BD",x"FC",x"A9",x"9D",x"24",x"19", -- 0x0500
    x"CA",x"10",x"F7",x"60",x"C6",x"7C",x"10",x"2E", -- 0x0508
    x"A9",x"0C",x"85",x"7C",x"A9",x"FB",x"8D",x"20", -- 0x0510
    x"91",x"AD",x"21",x"91",x"30",x"0B",x"AD",x"00", -- 0x0518
    x"90",x"18",x"69",x"01",x"29",x"8F",x"8D",x"00", -- 0x0520
    x"90",x"A9",x"F7",x"8D",x"20",x"91",x"AD",x"21", -- 0x0528
    x"91",x"30",x"0B",x"AD",x"01",x"90",x"18",x"69", -- 0x0530
    x"01",x"29",x"1F",x"8D",x"01",x"90",x"A5",x"8B", -- 0x0538
    x"F0",x"0B",x"20",x"80",x"A5",x"F0",x"34",x"A9", -- 0x0540
    x"00",x"85",x"8B",x"F0",x"2E",x"20",x"80",x"A5", -- 0x0548
    x"D0",x"0E",x"AD",x"00",x"90",x"49",x"80",x"8D", -- 0x0550
    x"00",x"90",x"A9",x"FF",x"85",x"8B",x"D0",x"1B", -- 0x0558
    x"A9",x"EF",x"8D",x"20",x"91",x"AD",x"21",x"91", -- 0x0560
    x"30",x"04",x"A9",x"01",x"D0",x"0F",x"A9",x"DF", -- 0x0568
    x"8D",x"20",x"91",x"AD",x"21",x"91",x"30",x"03", -- 0x0570
    x"A9",x"03",x"2C",x"A9",x"00",x"85",x"68",x"60", -- 0x0578
    x"A9",x"7F",x"8D",x"20",x"91",x"AD",x"21",x"91", -- 0x0580
    x"29",x"80",x"D0",x"16",x"A9",x"F7",x"8D",x"20", -- 0x0588
    x"91",x"AD",x"21",x"91",x"29",x"02",x"F0",x"0A", -- 0x0590
    x"A9",x"EF",x"8D",x"20",x"91",x"AD",x"21",x"91", -- 0x0598
    x"29",x"40",x"60",x"20",x"96",x"A8",x"20",x"0C", -- 0x05A0
    x"A5",x"A5",x"68",x"D0",x"F6",x"20",x"96",x"A8", -- 0x05A8
    x"20",x"0C",x"A5",x"A5",x"68",x"F0",x"F6",x"60", -- 0x05B0
    x"48",x"20",x"C0",x"A5",x"20",x"A8",x"A8",x"68", -- 0x05B8
    x"AA",x"D0",x"0B",x"A0",x"2B",x"B9",x"00",x"18", -- 0x05C0
    x"99",x"BF",x"00",x"88",x"10",x"F7",x"A9",x"93", -- 0x05C8
    x"20",x"2E",x"B2",x"A0",x"2B",x"B9",x"A0",x"A9", -- 0x05D0
    x"99",x"00",x"18",x"A9",x"03",x"99",x"00",x"94", -- 0x05D8
    x"88",x"10",x"F2",x"8A",x"D0",x"0A",x"A2",x"2B", -- 0x05E0
    x"B5",x"BF",x"9D",x"00",x"18",x"CA",x"10",x"F8", -- 0x05E8
    x"A0",x"01",x"A2",x"15",x"A9",x"52",x"20",x"AE", -- 0x05F0
    x"A7",x"A9",x"03",x"20",x"C4",x"A7",x"CA",x"10", -- 0x05F8
    x"F3",x"C8",x"A2",x"00",x"A9",x"50",x"20",x"AE", -- 0x0600
    x"A7",x"A9",x"03",x"20",x"C4",x"A7",x"A2",x"15", -- 0x0608
    x"A9",x"51",x"20",x"AE",x"A7",x"A9",x"03",x"20", -- 0x0610
    x"C4",x"A7",x"C8",x"C0",x"19",x"D0",x"E3",x"A2", -- 0x0618
    x"02",x"A9",x"5B",x"A0",x"10",x"20",x"AE",x"A7", -- 0x0620
    x"A9",x"03",x"20",x"C4",x"A7",x"A0",x"14",x"A9", -- 0x0628
    x"5B",x"20",x"AE",x"A7",x"A9",x"03",x"20",x"C4", -- 0x0630
    x"A7",x"CA",x"D0",x"E5",x"A2",x"13",x"A9",x"5B", -- 0x0638
    x"A0",x"10",x"20",x"AE",x"A7",x"A9",x"03",x"20", -- 0x0640
    x"C4",x"A7",x"A0",x"14",x"A9",x"5B",x"20",x"AE", -- 0x0648
    x"A7",x"A9",x"03",x"20",x"C4",x"A7",x"E8",x"E0", -- 0x0650
    x"15",x"D0",x"E3",x"A2",x"14",x"A9",x"06",x"9D", -- 0x0658
    x"58",x"94",x"A9",x"05",x"9D",x"84",x"94",x"A9", -- 0x0660
    x"07",x"9D",x"B0",x"94",x"CA",x"D0",x"EE",x"A0", -- 0x0668
    x"02",x"20",x"6C",x"A3",x"88",x"10",x"FA",x"A9", -- 0x0670
    x"09",x"85",x"98",x"85",x"99",x"85",x"9A",x"60", -- 0x0678
    x"85",x"96",x"98",x"48",x"8A",x"48",x"A5",x"96", -- 0x0680
    x"30",x"30",x"A2",x"09",x"A9",x"20",x"9D",x"92", -- 0x0688
    x"19",x"CA",x"10",x"FA",x"A5",x"96",x"29",x"40", -- 0x0690
    x"F0",x"0B",x"A2",x"09",x"BD",x"D2",x"A9",x"9D", -- 0x0698
    x"92",x"19",x"CA",x"10",x"F7",x"A5",x"96",x"29", -- 0x06A0
    x"01",x"18",x"69",x"31",x"8D",x"6E",x"19",x"A2", -- 0x06A8
    x"05",x"BD",x"CC",x"A9",x"9D",x"67",x"19",x"CA", -- 0x06B0
    x"10",x"F7",x"A2",x"1E",x"A9",x"00",x"95",x"73", -- 0x06B8
    x"CA",x"10",x"FB",x"68",x"C9",x"58",x"90",x"08", -- 0x06C0
    x"69",x"0B",x"A2",x"FF",x"A0",x"04",x"D0",x"06", -- 0x06C8
    x"E9",x"0B",x"A2",x"01",x"A0",x"06",x"48",x"86", -- 0x06D0
    x"89",x"84",x"7F",x"A9",x"0B",x"85",x"80",x"A9", -- 0x06D8
    x"0A",x"85",x"81",x"20",x"34",x"A2",x"A5",x"96", -- 0x06E0
    x"30",x"08",x"A6",x"95",x"20",x"8C",x"A1",x"4C", -- 0x06E8
    x"F5",x"A6",x"20",x"E5",x"A4",x"20",x"96",x"A8", -- 0x06F0
    x"C6",x"81",x"D0",x"E7",x"68",x"AA",x"68",x"48", -- 0x06F8
    x"A8",x"8A",x"48",x"20",x"4C",x"A0",x"A5",x"7F", -- 0x0700
    x"49",x"01",x"85",x"7F",x"68",x"18",x"65",x"89", -- 0x0708
    x"48",x"C6",x"80",x"D0",x"CA",x"A2",x"07",x"A9", -- 0x0710
    x"20",x"9D",x"67",x"19",x"CA",x"10",x"FA",x"68", -- 0x0718
    x"68",x"60",x"A9",x"02",x"85",x"74",x"A0",x"02", -- 0x0720
    x"A2",x"01",x"86",x"73",x"84",x"74",x"A9",x"20", -- 0x0728
    x"20",x"AE",x"A7",x"E8",x"E0",x"15",x"D0",x"F2", -- 0x0730
    x"C8",x"C0",x"19",x"D0",x"EB",x"A9",x"02",x"85", -- 0x0738
    x"74",x"A0",x"00",x"A2",x"00",x"A9",x"01",x"85", -- 0x0740
    x"73",x"B9",x"58",x"AC",x"85",x"72",x"B9",x"6D", -- 0x0748
    x"AC",x"85",x"76",x"BD",x"81",x"AB",x"30",x"16", -- 0x0750
    x"20",x"B2",x"A7",x"A5",x"73",x"C5",x"76",x"B0", -- 0x0758
    x"03",x"A5",x"72",x"2C",x"A9",x"01",x"20",x"C8", -- 0x0760
    x"A7",x"E6",x"73",x"E8",x"D0",x"E5",x"C9",x"FF", -- 0x0768
    x"F0",x"06",x"E8",x"C8",x"E6",x"74",x"D0",x"CD", -- 0x0770
    x"A0",x"05",x"A2",x"4E",x"20",x"0C",x"A5",x"C9", -- 0x0778
    x"01",x"F0",x"0E",x"20",x"96",x"A8",x"CA",x"D0", -- 0x0780
    x"F3",x"88",x"D0",x"F0",x"A9",x"00",x"85",x"68", -- 0x0788
    x"60",x"A9",x"FF",x"85",x"68",x"60",x"48",x"8A", -- 0x0790
    x"48",x"A6",x"74",x"BD",x"5E",x"A9",x"18",x"65", -- 0x0798
    x"73",x"85",x"6E",x"BD",x"79",x"A9",x"69",x"00", -- 0x07A0
    x"85",x"6F",x"68",x"AA",x"68",x"60",x"86",x"73", -- 0x07A8
    x"84",x"74",x"85",x"78",x"98",x"48",x"A5",x"78", -- 0x07B0
    x"20",x"96",x"A7",x"A0",x"00",x"91",x"6E",x"68", -- 0x07B8
    x"A8",x"A5",x"78",x"60",x"86",x"73",x"84",x"74", -- 0x07C0
    x"85",x"78",x"98",x"48",x"20",x"96",x"A7",x"A5", -- 0x07C8
    x"6F",x"18",x"69",x"7C",x"85",x"6F",x"A5",x"78", -- 0x07D0
    x"A0",x"00",x"91",x"6E",x"68",x"A8",x"A5",x"78", -- 0x07D8
    x"60",x"85",x"72",x"A9",x"01",x"85",x"7B",x"98", -- 0x07E0
    x"48",x"30",x"03",x"A9",x"00",x"2C",x"A9",x"0F", -- 0x07E8
    x"85",x"7A",x"A5",x"72",x"20",x"1A",x"A8",x"A2", -- 0x07F0
    x"0A",x"A0",x"00",x"68",x"29",x"7F",x"09",x"70", -- 0x07F8
    x"4C",x"AE",x"A7",x"48",x"8A",x"48",x"A2",x"00", -- 0x0800
    x"BD",x"F2",x"A9",x"20",x"2E",x"B2",x"E8",x"E0", -- 0x0808
    x"0A",x"D0",x"F5",x"68",x"AA",x"68",x"A0",x"00", -- 0x0810
    x"84",x"7B",x"A0",x"00",x"84",x"79",x"A0",x"05", -- 0x0818
    x"48",x"A9",x"00",x"85",x"72",x"68",x"38",x"F9", -- 0x0820
    x"64",x"A8",x"48",x"8A",x"F9",x"69",x"A8",x"AA", -- 0x0828
    x"68",x"90",x"04",x"E6",x"72",x"D0",x"EF",x"79", -- 0x0830
    x"64",x"A8",x"48",x"8A",x"79",x"69",x"A8",x"AA", -- 0x0838
    x"68",x"E6",x"72",x"C6",x"72",x"D0",x"0F",x"E6", -- 0x0840
    x"79",x"C6",x"79",x"D0",x"09",x"C0",x"00",x"F0", -- 0x0848
    x"05",x"48",x"A9",x"20",x"D0",x"07",x"48",x"A5", -- 0x0850
    x"72",x"09",x"30",x"E6",x"79",x"20",x"6F",x"A8", -- 0x0858
    x"68",x"88",x"10",x"BC",x"60",x"01",x"0A",x"64", -- 0x0860
    x"E8",x"10",x"00",x"00",x"00",x"03",x"27",x"85", -- 0x0868
    x"78",x"8A",x"48",x"A5",x"78",x"A6",x"7B",x"D0", -- 0x0870
    x"06",x"20",x"2E",x"B2",x"4C",x"91",x"A8",x"A6", -- 0x0878
    x"7A",x"E6",x"7A",x"C9",x"20",x"D0",x"05",x"A9", -- 0x0880
    x"5F",x"4C",x"8E",x"A8",x"09",x"40",x"9D",x"16", -- 0x0888
    x"18",x"68",x"AA",x"A5",x"78",x"60",x"AD",x"1D", -- 0x0890
    x"91",x"29",x"40",x"F0",x"F9",x"A9",x"10",x"8D", -- 0x0898
    x"14",x"91",x"A9",x"27",x"8D",x"15",x"91",x"60", -- 0x08A0
    x"A2",x"02",x"B5",x"98",x"48",x"BD",x"00",x"14", -- 0x08A8
    x"95",x"98",x"68",x"9D",x"00",x"14",x"CA",x"10", -- 0x08B0
    x"F1",x"A2",x"1D",x"B5",x"A1",x"48",x"BD",x"03", -- 0x08B8
    x"14",x"95",x"A1",x"68",x"9D",x"03",x"14",x"CA", -- 0x08C0
    x"10",x"F1",x"A2",x"13",x"A9",x"20",x"9D",x"61", -- 0x08C8
    x"19",x"CA",x"10",x"FA",x"60",x"78",x"D8",x"A2", -- 0x08D0
    x"FF",x"9A",x"20",x"8A",x"FF",x"D8",x"78",x"A9", -- 0x08D8
    x"00",x"8D",x"1E",x"91",x"A9",x"7F",x"8D",x"2E", -- 0x08E0
    x"91",x"A9",x"00",x"8D",x"1B",x"91",x"8D",x"2B", -- 0x08E8
    x"91",x"A9",x"FF",x"8D",x"22",x"91",x"A9",x"80", -- 0x08F0
    x"8D",x"13",x"91",x"A2",x"00",x"8E",x"14",x"91", -- 0x08F8
    x"E8",x"8E",x"15",x"91",x"AD",x"1C",x"91",x"29", -- 0x0900
    x"3F",x"8D",x"1C",x"91",x"A2",x"0F",x"BD",x"4E", -- 0x0908
    x"A9",x"9D",x"00",x"90",x"CA",x"10",x"F7",x"A2", -- 0x0910
    x"00",x"8A",x"95",x"00",x"9D",x"00",x"1C",x"CA", -- 0x0918
    x"D0",x"F8",x"A2",x"00",x"BD",x"82",x"AC",x"9D", -- 0x0920
    x"00",x"10",x"BD",x"82",x"AD",x"9D",x"00",x"11", -- 0x0928
    x"BD",x"82",x"AE",x"9D",x"80",x"12",x"CA",x"D0", -- 0x0930
    x"EB",x"A9",x"FF",x"8D",x"80",x"13",x"BD",x"80", -- 0x0938
    x"11",x"49",x"FF",x"9D",x"81",x"13",x"E8",x"E0", -- 0x0940
    x"50",x"D0",x"F3",x"4C",x"00",x"B0",x"03",x"16", -- 0x0948
    x"16",x"34",x"00",x"EC",x"00",x"00",x"00",x"00", -- 0x0950
    x"00",x"00",x"00",x"00",x"00",x"0B",x"16",x"2C", -- 0x0958
    x"42",x"58",x"6E",x"84",x"9A",x"B0",x"C6",x"DC", -- 0x0960
    x"F2",x"08",x"1E",x"34",x"4A",x"60",x"76",x"8C", -- 0x0968
    x"A2",x"B8",x"CE",x"E4",x"FA",x"10",x"26",x"3C", -- 0x0970
    x"52",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0978
    x"18",x"18",x"18",x"18",x"19",x"19",x"19",x"19", -- 0x0980
    x"19",x"19",x"19",x"19",x"19",x"19",x"19",x"19", -- 0x0988
    x"1A",x"1A",x"1A",x"1A",x"00",x"16",x"2C",x"01", -- 0x0990
    x"17",x"2D",x"00",x"0A",x"14",x"0A",x"05",x"02", -- 0x0998
    x"21",x"22",x"23",x"24",x"25",x"26",x"71",x"5F", -- 0x09A0
    x"1B",x"1C",x"1D",x"21",x"1E",x"5F",x"5F",x"21", -- 0x09A8
    x"22",x"23",x"24",x"25",x"26",x"72",x"5F",x"5F", -- 0x09B0
    x"5F",x"5F",x"5F",x"70",x"5F",x"5F",x"5F",x"5F", -- 0x09B8
    x"70",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F", -- 0x09C0
    x"5F",x"5F",x"5F",x"5F",x"10",x"0C",x"01",x"19", -- 0x09C8
    x"05",x"12",x"02",x"0F",x"0E",x"15",x"13",x"20", -- 0x09D0
    x"10",x"0C",x"01",x"19",x"02",x"0F",x"0E",x"15", -- 0x09D8
    x"13",x"20",x"0A",x"15",x"0D",x"10",x"31",x"30", -- 0x09E0
    x"30",x"30",x"30",x"35",x"30",x"30",x"30",x"32", -- 0x09E8
    x"30",x"30",x"48",x"49",x"47",x"48",x"20",x"53", -- 0x09F0
    x"43",x"4F",x"52",x"45",x"07",x"01",x"0D",x"05", -- 0x09F8
    x"20",x"0F",x"16",x"05",x"12",x"E4",x"36",x"E4", -- 0x0A00
    x"12",x"E4",x"7E",x"E4",x"12",x"E7",x"12",x"E4", -- 0x0A08
    x"12",x"E7",x"12",x"EA",x"A2",x"00",x"E1",x"12", -- 0x0A10
    x"DF",x"12",x"E1",x"12",x"E8",x"24",x"E1",x"12", -- 0x0A18
    x"DB",x"24",x"DB",x"12",x"D9",x"12",x"DB",x"12", -- 0x0A20
    x"E1",x"24",x"DB",x"12",x"D2",x"24",x"DB",x"12", -- 0x0A28
    x"D7",x"12",x"D2",x"12",x"D7",x"24",x"D7",x"12", -- 0x0A30
    x"D7",x"24",x"DD",x"12",x"DB",x"12",x"D7",x"12", -- 0x0A38
    x"E1",x"24",x"DB",x"12",x"D2",x"24",x"00",x"BF", -- 0x0A40
    x"24",x"BF",x"18",x"BF",x"0C",x"BF",x"24",x"C9", -- 0x0A48
    x"20",x"C6",x"0C",x"C6",x"18",x"BF",x"0C",x"BF", -- 0x0A50
    x"18",x"BB",x"0C",x"BF",x"30",x"00",x"00",x"11", -- 0x0A58
    x"42",x"10",x"38",x"38",x"10",x"7C",x"BA",x"BA", -- 0x0A60
    x"BA",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A68
    x"00",x"7C",x"38",x"28",x"28",x"28",x"28",x"2F", -- 0x0A70
    x"F0",x"00",x"00",x"00",x"00",x"0F",x"F1",x"01", -- 0x0A78
    x"03",x"00",x"00",x"0F",x"F0",x"80",x"80",x"80", -- 0x0A80
    x"C0",x"0F",x"F0",x"00",x"00",x"00",x"00",x"00", -- 0x0A88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A90
    x"00",x"08",x"1C",x"1C",x"08",x"3E",x"5D",x"5D", -- 0x0A98
    x"5D",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AA0
    x"00",x"F0",x"0F",x"00",x"00",x"00",x"00",x"00", -- 0x0AA8
    x"00",x"00",x"00",x"F0",x"0F",x"01",x"01",x"01", -- 0x0AB0
    x"03",x"00",x"00",x"00",x"00",x"F0",x"8F",x"80", -- 0x0AB8
    x"C0",x"3E",x"1C",x"14",x"14",x"14",x"14",x"F4", -- 0x0AC0
    x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AC8
    x"00",x"92",x"BA",x"BA",x"54",x"7C",x"38",x"38", -- 0x0AD0
    x"38",x"38",x"38",x"44",x"44",x"82",x"82",x"82", -- 0x0AD8
    x"82",x"90",x"B8",x"B8",x"50",x"7C",x"3C",x"3A", -- 0x0AE0
    x"3A",x"3A",x"38",x"48",x"48",x"88",x"84",x"84", -- 0x0AE8
    x"84",x"10",x"38",x"38",x"10",x"7C",x"7C",x"BA", -- 0x0AF0
    x"BA",x"BA",x"38",x"28",x"28",x"28",x"44",x"44", -- 0x0AF8
    x"44",x"12",x"3A",x"3A",x"14",x"7C",x"78",x"B8", -- 0x0B00
    x"B8",x"B8",x"38",x"24",x"24",x"22",x"42",x"42", -- 0x0B08
    x"42",x"10",x"B8",x"B8",x"90",x"7C",x"3A",x"3A", -- 0x0B10
    x"3A",x"38",x"38",x"28",x"28",x"50",x"50",x"48", -- 0x0B18
    x"44",x"10",x"38",x"38",x"96",x"BA",x"FA",x"BA", -- 0x0B20
    x"38",x"38",x"38",x"28",x"48",x"90",x"90",x"8C", -- 0x0B28
    x"82",x"10",x"3A",x"3A",x"12",x"7C",x"B8",x"B8", -- 0x0B30
    x"B8",x"38",x"38",x"28",x"28",x"14",x"14",x"24", -- 0x0B38
    x"44",x"10",x"38",x"3A",x"D2",x"BA",x"BE",x"BA", -- 0x0B40
    x"38",x"38",x"38",x"28",x"24",x"12",x"12",x"62", -- 0x0B48
    x"82",x"92",x"BA",x"BA",x"54",x"7C",x"38",x"38", -- 0x0B50
    x"38",x"38",x"38",x"28",x"28",x"28",x"28",x"28", -- 0x0B58
    x"28",x"00",x"00",x"10",x"38",x"38",x"10",x"78", -- 0x0B60
    x"B8",x"B8",x"B8",x"B8",x"38",x"28",x"28",x"14", -- 0x0B68
    x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B70
    x"00",x"00",x"00",x"00",x"00",x"6E",x"FE",x"6F", -- 0x0B78
    x"09",x"80",x"20",x"20",x"20",x"09",x"0E",x"13", -- 0x0B80
    x"14",x"12",x"15",x"03",x"14",x"09",x"0F",x"0E", -- 0x0B88
    x"13",x"3A",x"80",x"80",x"80",x"13",x"03",x"0F", -- 0x0B90
    x"12",x"05",x"20",x"01",x"04",x"16",x"01",x"0E", -- 0x0B98
    x"03",x"05",x"20",x"20",x"14",x"01",x"02",x"0C", -- 0x0BA0
    x"05",x"80",x"80",x"20",x"20",x"20",x"20",x"0A", -- 0x0BA8
    x"15",x"0D",x"10",x"13",x"20",x"2D",x"20",x"31", -- 0x0BB0
    x"30",x"80",x"80",x"20",x"02",x"01",x"0C",x"0C", -- 0x0BB8
    x"0F",x"0F",x"0E",x"13",x"20",x"20",x"20",x"02", -- 0x0BC0
    x"0F",x"0E",x"15",x"13",x"80",x"80",x"20",x"20", -- 0x0BC8
    x"60",x"20",x"2D",x"20",x"32",x"30",x"20",x"20", -- 0x0BD0
    x"20",x"20",x"20",x"32",x"30",x"30",x"80",x"20", -- 0x0BD8
    x"20",x"60",x"20",x"2D",x"20",x"35",x"30",x"20", -- 0x0BE0
    x"20",x"20",x"20",x"20",x"35",x"30",x"30",x"80", -- 0x0BE8
    x"20",x"20",x"60",x"20",x"2D",x"31",x"30",x"30", -- 0x0BF0
    x"20",x"20",x"20",x"20",x"31",x"30",x"30",x"30", -- 0x0BF8
    x"2B",x"80",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x0C00
    x"20",x"20",x"20",x"02",x"0F",x"0E",x"15",x"13", -- 0x0C08
    x"20",x"0A",x"15",x"0D",x"10",x"80",x"28",x"0F", -- 0x0C10
    x"0E",x"03",x"05",x"20",x"06",x"0F",x"12",x"20", -- 0x0C18
    x"05",x"01",x"03",x"08",x"20",x"0A",x"15",x"0D", -- 0x0C20
    x"10",x"29",x"80",x"80",x"80",x"20",x"35",x"20", -- 0x0C28
    x"0A",x"15",x"0D",x"10",x"13",x"20",x"10",x"05", -- 0x0C30
    x"12",x"20",x"10",x"0C",x"01",x"19",x"05",x"12", -- 0x0C38
    x"80",x"80",x"80",x"20",x"28",x"03",x"29",x"20", -- 0x0C40
    x"31",x"39",x"38",x"32",x"20",x"03",x"0F",x"0D", -- 0x0C48
    x"0D",x"0F",x"04",x"0F",x"12",x"05",x"80",x"FF", -- 0x0C50
    x"00",x"01",x"00",x"00",x"03",x"00",x"07",x"00", -- 0x0C58
    x"01",x"00",x"07",x"05",x"06",x"01",x"01",x"00", -- 0x0C60
    x"00",x"05",x"00",x"00",x"03",x"00",x"16",x"00", -- 0x0C68
    x"00",x"16",x"00",x"16",x"00",x"16",x"00",x"05", -- 0x0C70
    x"05",x"05",x"16",x"16",x"00",x"00",x"16",x"00", -- 0x0C78
    x"00",x"16",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C80
    x"00",x"00",x"38",x"6C",x"C6",x"C6",x"FE",x"C6", -- 0x0C88
    x"C6",x"00",x"FC",x"66",x"66",x"7C",x"66",x"66", -- 0x0C90
    x"FC",x"00",x"3C",x"66",x"C0",x"C0",x"C0",x"66", -- 0x0C98
    x"3C",x"00",x"F8",x"64",x"66",x"66",x"66",x"64", -- 0x0CA0
    x"F8",x"00",x"FE",x"60",x"60",x"7C",x"60",x"60", -- 0x0CA8
    x"FE",x"00",x"FE",x"60",x"60",x"7C",x"60",x"60", -- 0x0CB0
    x"F0",x"00",x"3C",x"66",x"C0",x"DE",x"C6",x"66", -- 0x0CB8
    x"3C",x"00",x"C6",x"C6",x"C6",x"FE",x"C6",x"C6", -- 0x0CC0
    x"C6",x"00",x"3C",x"18",x"18",x"18",x"18",x"18", -- 0x0CC8
    x"3C",x"00",x"1E",x"0C",x"0C",x"0C",x"CC",x"CC", -- 0x0CD0
    x"78",x"00",x"C6",x"CC",x"D8",x"F0",x"D8",x"CC", -- 0x0CD8
    x"C6",x"00",x"F0",x"60",x"60",x"60",x"60",x"60", -- 0x0CE0
    x"FE",x"00",x"C6",x"EE",x"FE",x"D6",x"C6",x"C6", -- 0x0CE8
    x"C6",x"00",x"C6",x"E6",x"F6",x"DE",x"CE",x"C6", -- 0x0CF0
    x"C6",x"00",x"7C",x"EE",x"C6",x"C6",x"C6",x"EE", -- 0x0CF8
    x"7C",x"00",x"FC",x"66",x"66",x"7C",x"60",x"60", -- 0x0D00
    x"F0",x"00",x"38",x"64",x"C2",x"C2",x"CA",x"64", -- 0x0D08
    x"3A",x"00",x"FC",x"C6",x"C6",x"FC",x"D8",x"CC", -- 0x0D10
    x"C6",x"00",x"7C",x"C6",x"C0",x"7C",x"06",x"C6", -- 0x0D18
    x"7C",x"00",x"7E",x"18",x"18",x"18",x"18",x"18", -- 0x0D20
    x"3C",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6", -- 0x0D28
    x"7C",x"00",x"C6",x"C6",x"C6",x"6C",x"6C",x"38", -- 0x0D30
    x"38",x"00",x"C6",x"C6",x"C6",x"D6",x"D6",x"FE", -- 0x0D38
    x"6C",x"00",x"C6",x"C6",x"6C",x"38",x"6C",x"C6", -- 0x0D40
    x"C6",x"00",x"C6",x"C6",x"6C",x"7C",x"38",x"38", -- 0x0D48
    x"38",x"00",x"FE",x"C6",x"0C",x"38",x"60",x"C6", -- 0x0D50
    x"FE",x"00",x"FF",x"E1",x"F3",x"F3",x"F3",x"33", -- 0x0D58
    x"33",x"87",x"FF",x"39",x"39",x"39",x"39",x"39", -- 0x0D60
    x"39",x"83",x"FF",x"39",x"11",x"01",x"29",x"39", -- 0x0D68
    x"39",x"39",x"FF",x"83",x"39",x"3F",x"83",x"F9", -- 0x0D70
    x"39",x"83",x"00",x"20",x"40",x"FE",x"FE",x"40", -- 0x0D78
    x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D80
    x"00",x"00",x"FF",x"03",x"99",x"99",x"83",x"9F", -- 0x0D88
    x"9F",x"0F",x"FF",x"0F",x"9F",x"9F",x"9F",x"9F", -- 0x0D90
    x"9F",x"01",x"FF",x"C7",x"93",x"39",x"39",x"01", -- 0x0D98
    x"39",x"39",x"FF",x"39",x"39",x"93",x"83",x"C7", -- 0x0DA0
    x"C7",x"C7",x"FF",x"01",x"9F",x"9F",x"83",x"9F", -- 0x0DA8
    x"9F",x"01",x"FF",x"03",x"39",x"39",x"03",x"27", -- 0x0DB0
    x"33",x"39",x"0C",x"18",x"30",x"00",x"00",x"00", -- 0x0DB8
    x"00",x"00",x"0C",x"18",x"30",x"30",x"30",x"18", -- 0x0DC0
    x"0C",x"00",x"30",x"18",x"0C",x"0C",x"0C",x"18", -- 0x0DC8
    x"30",x"00",x"10",x"54",x"38",x"FE",x"38",x"54", -- 0x0DD0
    x"10",x"00",x"00",x"18",x"18",x"7E",x"7E",x"18", -- 0x0DD8
    x"18",x"00",x"00",x"00",x"00",x"00",x"18",x"18", -- 0x0DE0
    x"30",x"60",x"00",x"00",x"00",x"7E",x"7E",x"00", -- 0x0DE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- 0x0DF0
    x"18",x"00",x"00",x"06",x"0C",x"18",x"30",x"60", -- 0x0DF8
    x"C0",x"00",x"7C",x"C6",x"CE",x"D6",x"E6",x"C6", -- 0x0E00
    x"7C",x"00",x"18",x"38",x"18",x"18",x"18",x"18", -- 0x0E08
    x"3C",x"00",x"7C",x"C6",x"C6",x"0C",x"38",x"E0", -- 0x0E10
    x"FE",x"00",x"7C",x"C6",x"06",x"1C",x"06",x"C6", -- 0x0E18
    x"7C",x"00",x"0C",x"1C",x"2C",x"4C",x"FE",x"0C", -- 0x0E20
    x"0C",x"00",x"FE",x"C0",x"C0",x"FC",x"06",x"C6", -- 0x0E28
    x"7C",x"00",x"1C",x"30",x"60",x"FC",x"C6",x"C6", -- 0x0E30
    x"7C",x"00",x"7E",x"C6",x"0C",x"18",x"18",x"18", -- 0x0E38
    x"18",x"00",x"7C",x"C6",x"C6",x"7C",x"C6",x"C6", -- 0x0E40
    x"7C",x"00",x"7C",x"C6",x"C6",x"7E",x"06",x"0C", -- 0x0E48
    x"38",x"00",x"00",x"18",x"18",x"00",x"18",x"18", -- 0x0E50
    x"00",x"00",x"00",x"18",x"18",x"00",x"18",x"18", -- 0x0E58
    x"20",x"00",x"06",x"0C",x"18",x"30",x"18",x"0C", -- 0x0E60
    x"06",x"00",x"00",x"00",x"7E",x"00",x"7E",x"00", -- 0x0E68
    x"00",x"00",x"C0",x"60",x"30",x"18",x"30",x"60", -- 0x0E70
    x"C0",x"00",x"7C",x"C6",x"0C",x"18",x"00",x"18", -- 0x0E78
    x"18",x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE", -- 0x0E80
    x"FE",x"FE",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F", -- 0x0E88
    x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E98
    x"FF",x"FF",x"30",x"30",x"A9",x"00",x"8D",x"22", -- 0x0EA0
    x"91",x"AD",x"20",x"91",x"2A",x"B0",x"09",x"A5", -- 0x0EA8
    x"FF",x"38",x"E9",x"03",x"90",x"02",x"85",x"FF", -- 0x0EB0
    x"AD",x"11",x"91",x"29",x"10",x"C9",x"10",x"F0", -- 0x0EB8
    x"09",x"A5",x"FF",x"18",x"69",x"03",x"B0",x"02", -- 0x0EC0
    x"85",x"FF",x"A9",x"FF",x"8D",x"22",x"91",x"A5", -- 0x0EC8
    x"FF",x"60",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x0ED0
    x"AA",x"AA",x"FF",x"FF",x"00",x"00",x"00",x"00", -- 0x0ED8
    x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00", -- 0x0EE0
    x"00",x"00",x"FF",x"24",x"24",x"24",x"24",x"24", -- 0x0EE8
    x"04",x"8C",x"FF",x"3F",x"9F",x"9F",x"3F",x"FF", -- 0x0EF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EF8
    x"FF",x"FF",x"3C",x"7E",x"FF",x"FF",x"DF",x"66", -- 0x0F00
    x"3C",x"18",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F08
    x"00",x"00",x"1F",x"3F",x"7F",x"7F",x"6F",x"33", -- 0x0F10
    x"1E",x"0C",x"00",x"00",x"80",x"80",x"80",x"00", -- 0x0F18
    x"00",x"00",x"0F",x"1F",x"3F",x"3F",x"37",x"19", -- 0x0F20
    x"0F",x"06",x"00",x"80",x"C0",x"C0",x"C0",x"80", -- 0x0F28
    x"00",x"00",x"07",x"0F",x"1F",x"1F",x"1B",x"0C", -- 0x0F30
    x"07",x"03",x"80",x"C0",x"E0",x"E0",x"E0",x"C0", -- 0x0F38
    x"80",x"00",x"03",x"07",x"0F",x"0F",x"0D",x"06", -- 0x0F40
    x"03",x"01",x"C0",x"E0",x"F0",x"F0",x"F0",x"60", -- 0x0F48
    x"C0",x"80",x"01",x"03",x"07",x"07",x"06",x"03", -- 0x0F50
    x"01",x"00",x"E0",x"F0",x"F8",x"F8",x"F8",x"30", -- 0x0F58
    x"E0",x"C0",x"00",x"01",x"03",x"03",x"03",x"01", -- 0x0F60
    x"00",x"00",x"F0",x"F8",x"FC",x"FC",x"7C",x"98", -- 0x0F68
    x"F0",x"60",x"00",x"00",x"01",x"01",x"01",x"00", -- 0x0F70
    x"00",x"00",x"78",x"FC",x"FE",x"FE",x"BE",x"CC", -- 0x0F78
    x"78",x"30",x"52",x"32",x"31",x"17",x"4D",x"53", -- 0x0F80
    x"47",x"50",x"52",x"4E",x"31",x"0B",x"4D",x"55", -- 0x0F88
    x"4C",x"31",x"36",x"20",x"31",x"B7",x"4D",x"55", -- 0x0F90
    x"4C",x"31",x"36",x"41",x"31",x"BE",x"4D",x"55", -- 0x0F98
    x"4C",x"31",x"36",x"4C",x"31",x"C2",x"4D",x"55", -- 0x0FA0
    x"4C",x"31",x"36",x"53",x"31",x"D5",x"4D",x"55", -- 0x0FA8
    x"4C",x"41",x"53",x"31",x"07",x"24",x"4D",x"55", -- 0x0FB0
    x"4C",x"41",x"53",x"32",x"07",x"27",x"4D",x"55", -- 0x0FB8
    x"4C",x"41",x"53",x"4E",x"07",x"29",x"4D",x"55", -- 0x0FC0
    x"4C",x"4F",x"4F",x"50",x"30",x"71",x"4D",x"55", -- 0x0FC8
    x"4C",x"54",x"41",x"58",x"30",x"63",x"4E",x"45", -- 0x0FD0
    x"57",x"49",x"44",x"56",x"02",x"B4",x"4E",x"45", -- 0x0FD8
    x"57",x"49",x"54",x"4D",x"10",x"9D",x"4E",x"45", -- 0x0FE0
    x"57",x"4C",x"56",x"4C",x"10",x"A3",x"4E",x"4F", -- 0x0FE8
    x"41",x"52",x"47",x"20",x"0D",x"EC",x"4E",x"4F", -- 0x0FF0
    x"41",x"52",x"52",x"59",x"05",x"D7",x"4E",x"4F", -- 0x0FF8
    x"A9",x"00",x"A2",x"1C",x"85",x"01",x"86",x"02", -- 0x1000
    x"D8",x"4C",x"4A",x"B3",x"A5",x"01",x"91",x"01", -- 0x1008
    x"C8",x"A5",x"02",x"91",x"01",x"38",x"98",x"65", -- 0x1010
    x"01",x"85",x"01",x"90",x"02",x"E6",x"02",x"60", -- 0x1018
    x"48",x"38",x"A5",x"01",x"E9",x"02",x"85",x"01", -- 0x1020
    x"B0",x"02",x"C6",x"02",x"A0",x"01",x"B1",x"01", -- 0x1028
    x"AA",x"88",x"B1",x"01",x"85",x"01",x"86",x"02", -- 0x1030
    x"68",x"60",x"48",x"A5",x"65",x"A2",x"7D",x"20", -- 0x1038
    x"63",x"B0",x"18",x"69",x"01",x"90",x"01",x"E8", -- 0x1040
    x"85",x"65",x"8A",x"48",x"A5",x"66",x"A2",x"7D", -- 0x1048
    x"20",x"63",x"B0",x"85",x"60",x"68",x"18",x"65", -- 0x1050
    x"60",x"AA",x"85",x"66",x"68",x"20",x"63",x"B0", -- 0x1058
    x"E8",x"8A",x"60",x"85",x"60",x"8A",x"F0",x"19", -- 0x1060
    x"CA",x"86",x"61",x"A2",x"08",x"A9",x"00",x"66", -- 0x1068
    x"60",x"90",x"02",x"65",x"61",x"6A",x"66",x"60", -- 0x1070
    x"CA",x"D0",x"F6",x"85",x"5E",x"AA",x"A5",x"60", -- 0x1078
    x"60",x"85",x"5E",x"60",x"85",x"62",x"8A",x"D0", -- 0x1080
    x"05",x"86",x"62",x"AA",x"F0",x"1F",x"A2",x"00", -- 0x1088
    x"86",x"60",x"E8",x"0A",x"90",x"FC",x"85",x"61", -- 0x1090
    x"A5",x"62",x"66",x"61",x"C5",x"61",x"90",x"02", -- 0x1098
    x"E5",x"61",x"26",x"60",x"CA",x"D0",x"F3",x"85", -- 0x10A0
    x"5F",x"AA",x"A5",x"60",x"60",x"85",x"38",x"20", -- 0x10A8
    x"F5",x"B0",x"0D",x"45",x"52",x"52",x"20",x"44", -- 0x10B0
    x"49",x"56",x"30",x"00",x"4C",x"00",x"70",x"AA", -- 0x10B8
    x"A9",x"00",x"85",x"63",x"8A",x"A0",x"00",x"85", -- 0x10C0
    x"62",x"A5",x"5F",x"48",x"A2",x"0A",x"20",x"86", -- 0x10C8
    x"B0",x"85",x"62",x"8A",x"48",x"C8",x"A5",x"62", -- 0x10D0
    x"D0",x"F2",x"A5",x"63",x"F0",x"0A",x"84",x"63", -- 0x10D8
    x"38",x"E5",x"63",x"90",x"03",x"20",x"27",x"B1", -- 0x10E0
    x"68",x"09",x"30",x"20",x"33",x"B1",x"88",x"D0", -- 0x10E8
    x"F7",x"68",x"85",x"5F",x"60",x"68",x"85",x"34", -- 0x10F0
    x"68",x"85",x"35",x"20",x"0B",x"B1",x"38",x"98", -- 0x10F8
    x"65",x"34",x"85",x"34",x"90",x"02",x"E6",x"35", -- 0x1100
    x"6C",x"34",x"00",x"A0",x"01",x"B1",x"34",x"F0", -- 0x1108
    x"06",x"20",x"33",x"B1",x"C8",x"D0",x"F6",x"60", -- 0x1110
    x"A9",x"0D",x"4C",x"33",x"B1",x"AA",x"F0",x"F7", -- 0x1118
    x"20",x"18",x"B1",x"CA",x"D0",x"FA",x"60",x"AA", -- 0x1120
    x"F0",x"ED",x"A9",x"20",x"20",x"33",x"B1",x"CA", -- 0x1128
    x"D0",x"FA",x"60",x"85",x"63",x"48",x"8A",x"48", -- 0x1130
    x"98",x"48",x"A6",x"38",x"A0",x"00",x"20",x"47", -- 0x1138
    x"B1",x"68",x"A8",x"68",x"AA",x"68",x"60",x"E8", -- 0x1140
    x"CA",x"F0",x"04",x"C8",x"C8",x"D0",x"F9",x"B9", -- 0x1148
    x"86",x"B1",x"BE",x"87",x"B1",x"85",x"36",x"86", -- 0x1150
    x"37",x"A5",x"63",x"6C",x"36",x"00",x"20",x"0C", -- 0x1158
    x"B0",x"A0",x"00",x"B1",x"01",x"85",x"35",x"C8", -- 0x1160
    x"B1",x"01",x"85",x"34",x"C8",x"B1",x"01",x"85", -- 0x1168
    x"60",x"C8",x"B1",x"01",x"AA",x"C8",x"B1",x"01", -- 0x1170
    x"A8",x"A5",x"60",x"08",x"20",x"08",x"B1",x"28", -- 0x1178
    x"4C",x"20",x"B0",x"4C",x"D2",x"FF",x"83",x"B1", -- 0x1180
    x"2E",x"B2",x"83",x"B1",x"83",x"B1",x"83",x"B1", -- 0x1188
    x"83",x"B1",x"83",x"B1",x"83",x"B1",x"83",x"B1", -- 0x1190
    x"83",x"B1",x"20",x"0C",x"B0",x"A0",x"00",x"84", -- 0x1198
    x"5F",x"84",x"5E",x"B1",x"01",x"85",x"61",x"C8", -- 0x11A0
    x"B1",x"01",x"85",x"60",x"C8",x"B1",x"01",x"85", -- 0x11A8
    x"35",x"C8",x"B1",x"01",x"85",x"34",x"60",x"20", -- 0x11B0
    x"9A",x"B1",x"A2",x"10",x"D0",x"04",x"06",x"62", -- 0x11B8
    x"26",x"5E",x"06",x"60",x"26",x"61",x"90",x"0D", -- 0x11C0
    x"18",x"A5",x"34",x"65",x"62",x"85",x"62",x"A5", -- 0x11C8
    x"35",x"65",x"5E",x"85",x"5E",x"CA",x"D0",x"E6", -- 0x11D0
    x"A5",x"62",x"4C",x"20",x"B0",x"20",x"AD",x"B0", -- 0x11D8
    x"20",x"9A",x"B1",x"05",x"35",x"F0",x"F6",x"A5", -- 0x11E0
    x"60",x"05",x"61",x"F0",x"38",x"A2",x"11",x"CA", -- 0x11E8
    x"06",x"60",x"26",x"61",x"90",x"F9",x"26",x"62", -- 0x11F0
    x"26",x"5E",x"A5",x"62",x"C5",x"34",x"A5",x"5E", -- 0x11F8
    x"E5",x"35",x"90",x"09",x"85",x"5E",x"A5",x"62", -- 0x1200
    x"E5",x"34",x"85",x"62",x"38",x"26",x"60",x"26", -- 0x1208
    x"61",x"CA",x"D0",x"E2",x"A5",x"5E",x"85",x"64", -- 0x1210
    x"A5",x"62",x"85",x"5F",x"A5",x"61",x"85",x"5E", -- 0x1218
    x"A5",x"60",x"4C",x"20",x"B0",x"85",x"64",x"85", -- 0x1220
    x"5F",x"F0",x"F3",x"A5",x"64",x"60",x"48",x"85", -- 0x1228
    x"06",x"8A",x"48",x"98",x"48",x"A2",x"06",x"A5", -- 0x1230
    x"06",x"DD",x"80",x"B2",x"F0",x"36",x"CA",x"10", -- 0x1238
    x"F8",x"20",x"1E",x"B3",x"20",x"DB",x"B2",x"A5", -- 0x1240
    x"06",x"91",x"04",x"A5",x"05",x"18",x"69",x"7C", -- 0x1248
    x"85",x"05",x"A5",x"03",x"91",x"04",x"E6",x"07", -- 0x1250
    x"A5",x"07",x"C9",x"16",x"D0",x"10",x"A9",x"00", -- 0x1258
    x"85",x"07",x"E6",x"08",x"A5",x"08",x"C9",x"19", -- 0x1260
    x"D0",x"04",x"A9",x"00",x"85",x"08",x"68",x"A8", -- 0x1268
    x"68",x"AA",x"68",x"60",x"8A",x"0A",x"AA",x"BD", -- 0x1270
    x"88",x"B2",x"48",x"BD",x"87",x"B2",x"48",x"60", -- 0x1278
    x"9D",x"1D",x"91",x"11",x"13",x"0D",x"93",x"94", -- 0x1280
    x"B2",x"55",x"B2",x"9C",x"B2",x"61",x"B2",x"A6", -- 0x1288
    x"B2",x"AE",x"B2",x"B4",x"B2",x"C6",x"07",x"10", -- 0x1290
    x"D5",x"A9",x"15",x"85",x"07",x"C6",x"08",x"10", -- 0x1298
    x"CD",x"A9",x"18",x"85",x"08",x"D0",x"C7",x"A9", -- 0x12A0
    x"00",x"85",x"07",x"85",x"08",x"F0",x"BF",x"A9", -- 0x12A8
    x"00",x"85",x"07",x"F0",x"AD",x"A2",x"00",x"A9", -- 0x12B0
    x"20",x"9D",x"00",x"18",x"9D",x"00",x"19",x"9D", -- 0x12B8
    x"00",x"1A",x"9D",x"00",x"1B",x"E8",x"D0",x"F1", -- 0x12C0
    x"A9",x"01",x"9D",x"00",x"94",x"9D",x"00",x"95", -- 0x12C8
    x"9D",x"00",x"96",x"9D",x"00",x"97",x"E8",x"D0", -- 0x12D0
    x"F1",x"F0",x"CC",x"A5",x"08",x"0A",x"AA",x"BD", -- 0x12D8
    x"EC",x"B2",x"85",x"04",x"BD",x"ED",x"B2",x"85", -- 0x12E0
    x"05",x"A4",x"07",x"60",x"00",x"18",x"16",x"18", -- 0x12E8
    x"2C",x"18",x"42",x"18",x"58",x"18",x"6E",x"18", -- 0x12F0
    x"84",x"18",x"9A",x"18",x"B0",x"18",x"C6",x"18", -- 0x12F8
    x"DC",x"18",x"F2",x"18",x"08",x"19",x"1E",x"19", -- 0x1300
    x"34",x"19",x"4A",x"19",x"60",x"19",x"76",x"19", -- 0x1308
    x"8C",x"19",x"A2",x"19",x"B8",x"19",x"CE",x"19", -- 0x1310
    x"E4",x"19",x"FA",x"19",x"10",x"1A",x"A5",x"06", -- 0x1318
    x"30",x"05",x"29",x"3F",x"85",x"06",x"60",x"29", -- 0x1320
    x"3F",x"09",x"40",x"D0",x"F7",x"20",x"0C",x"B0", -- 0x1328
    x"A0",x"00",x"B1",x"01",x"85",x"07",x"C8",x"B1", -- 0x1330
    x"01",x"85",x"08",x"4C",x"20",x"B0",x"20",x"0C", -- 0x1338
    x"B0",x"A0",x"00",x"B1",x"01",x"85",x"03",x"4C", -- 0x1340
    x"20",x"B0",x"A0",x"43",x"20",x"44",x"B4",x"A0", -- 0x1348
    x"43",x"20",x"6C",x"BC",x"A0",x"43",x"20",x"87", -- 0x1350
    x"BE",x"A9",x"FF",x"8D",x"12",x"1C",x"A9",x"18", -- 0x1358
    x"A0",x"45",x"91",x"01",x"A0",x"43",x"20",x"BA", -- 0x1360
    x"BA",x"A9",x"00",x"8D",x"1D",x"1C",x"8D",x"1F", -- 0x1368
    x"1C",x"8D",x"1C",x"1C",x"8D",x"1E",x"1C",x"A0", -- 0x1370
    x"43",x"20",x"E6",x"B4",x"A0",x"43",x"20",x"76", -- 0x1378
    x"B5",x"A0",x"43",x"20",x"18",x"BB",x"AD",x"20", -- 0x1380
    x"1C",x"0D",x"21",x"1C",x"C9",x"00",x"F0",x"04", -- 0x1388
    x"A9",x"00",x"F0",x"02",x"A9",x"FF",x"F0",x"E4", -- 0x1390
    x"A9",x"06",x"A0",x"45",x"91",x"01",x"A9",x"10", -- 0x1398
    x"C8",x"91",x"01",x"A0",x"43",x"20",x"2D",x"B3", -- 0x13A0
    x"A9",x"01",x"85",x"38",x"20",x"F5",x"B0",x"47", -- 0x13A8
    x"41",x"4D",x"45",x"20",x"4F",x"56",x"45",x"52", -- 0x13B0
    x"00",x"A9",x"FF",x"A0",x"45",x"91",x"01",x"A0", -- 0x13B8
    x"43",x"20",x"5B",x"BE",x"A9",x"00",x"8D",x"13", -- 0x13C0
    x"1C",x"A9",x"01",x"48",x"AD",x"13",x"1C",x"A8", -- 0x13C8
    x"B9",x"1C",x"1C",x"18",x"ED",x"10",x"1C",x"B0", -- 0x13D0
    x"04",x"A9",x"00",x"F0",x"02",x"A9",x"FF",x"48", -- 0x13D8
    x"AD",x"13",x"1C",x"A8",x"B9",x"1C",x"1C",x"CD", -- 0x13E0
    x"10",x"1C",x"F0",x"04",x"A9",x"00",x"F0",x"02", -- 0x13E8
    x"A9",x"FF",x"48",x"AD",x"13",x"1C",x"A8",x"B9", -- 0x13F0
    x"1E",x"1C",x"18",x"ED",x"11",x"1C",x"B0",x"04", -- 0x13F8
    x"A9",x"00",x"F0",x"02",x"A9",x"FF",x"85",x"60", -- 0x1400
    x"68",x"25",x"60",x"85",x"60",x"68",x"05",x"60", -- 0x1408
    x"D0",x"03",x"4C",x"29",x"B4",x"AD",x"13",x"1C", -- 0x1410
    x"A8",x"B9",x"1C",x"1C",x"8D",x"10",x"1C",x"AD", -- 0x1418
    x"13",x"1C",x"A8",x"B9",x"1E",x"1C",x"8D",x"11", -- 0x1420
    x"1C",x"BA",x"E8",x"AD",x"13",x"1C",x"DD",x"00", -- 0x1428
    x"01",x"B0",x"06",x"EE",x"13",x"1C",x"4C",x"CC", -- 0x1430
    x"B3",x"9A",x"A9",x"00",x"D0",x"03",x"4C",x"4F", -- 0x1438
    x"B3",x"4C",x"00",x"70",x"20",x"0C",x"B0",x"A9", -- 0x1440
    x"40",x"8D",x"2C",x"1C",x"A9",x"01",x"8D",x"28", -- 0x1448
    x"1C",x"A9",x"00",x"8D",x"34",x"1C",x"A9",x"06", -- 0x1450
    x"8D",x"30",x"1C",x"A9",x"C0",x"8D",x"2D",x"1C", -- 0x1458
    x"A9",x"00",x"8D",x"29",x"1C",x"A9",x"60",x"8D", -- 0x1460
    x"35",x"1C",x"A9",x"06",x"8D",x"31",x"1C",x"A9", -- 0x1468
    x"E0",x"8D",x"2E",x"1C",x"A9",x"00",x"8D",x"2A", -- 0x1470
    x"1C",x"A9",x"28",x"8D",x"36",x"1C",x"A9",x"06", -- 0x1478
    x"8D",x"32",x"1C",x"A9",x"00",x"8D",x"2F",x"1C", -- 0x1480
    x"A9",x"FF",x"8D",x"2B",x"1C",x"A9",x"80",x"8D", -- 0x1488
    x"37",x"1C",x"A9",x"05",x"8D",x"33",x"1C",x"A9", -- 0x1490
    x"03",x"8D",x"25",x"1C",x"A9",x"0B",x"8D",x"26", -- 0x1498
    x"1C",x"A9",x"1B",x"8D",x"27",x"1C",x"A9",x"05", -- 0x14A0
    x"8D",x"3B",x"1C",x"A9",x"0C",x"8D",x"3C",x"1C", -- 0x14A8
    x"A9",x"1E",x"8D",x"3D",x"1C",x"A9",x"01",x"8D", -- 0x14B0
    x"38",x"1C",x"A9",x"02",x"8D",x"39",x"1C",x"A9", -- 0x14B8
    x"01",x"8D",x"3A",x"1C",x"A9",x"64",x"8D",x"40", -- 0x14C0
    x"1C",x"A9",x"32",x"8D",x"41",x"1C",x"A9",x"14", -- 0x14C8
    x"8D",x"42",x"1C",x"A9",x"0A",x"A0",x"03",x"91", -- 0x14D0
    x"01",x"A9",x"FF",x"C8",x"91",x"01",x"A0",x"01", -- 0x14D8
    x"20",x"BA",x"BA",x"4C",x"20",x"B0",x"20",x"0C", -- 0x14E0
    x"B0",x"A9",x"0A",x"A0",x"02",x"91",x"01",x"AD", -- 0x14E8
    x"12",x"1C",x"C8",x"91",x"01",x"A0",x"00",x"20", -- 0x14F0
    x"BA",x"BA",x"AD",x"0F",x"1C",x"29",x"01",x"8D", -- 0x14F8
    x"0C",x"1C",x"A9",x"00",x"48",x"AD",x"0C",x"1C", -- 0x1500
    x"48",x"A9",x"05",x"AA",x"68",x"A8",x"8A",x"99", -- 0x1508
    x"20",x"1C",x"AD",x"0C",x"1C",x"48",x"A9",x"FF", -- 0x1510
    x"AA",x"68",x"A8",x"8A",x"99",x"3E",x"1C",x"A0", -- 0x1518
    x"00",x"20",x"26",x"BC",x"68",x"CD",x"0C",x"1C", -- 0x1520
    x"B0",x"07",x"48",x"CE",x"0C",x"1C",x"4C",x"05", -- 0x1528
    x"B5",x"A9",x"00",x"8D",x"0D",x"1C",x"A9",x"01", -- 0x1530
    x"A0",x"02",x"91",x"01",x"A0",x"00",x"20",x"3E", -- 0x1538
    x"B3",x"AD",x"12",x"1C",x"D0",x"03",x"4C",x"73", -- 0x1540
    x"B5",x"A9",x"12",x"A0",x"02",x"91",x"01",x"A9", -- 0x1548
    x"08",x"C8",x"91",x"01",x"A9",x"54",x"C8",x"91", -- 0x1550
    x"01",x"A9",x"96",x"C8",x"91",x"01",x"A0",x"00", -- 0x1558
    x"20",x"BA",x"BA",x"A9",x"13",x"A0",x"02",x"91", -- 0x1560
    x"01",x"A9",x"00",x"C8",x"91",x"01",x"A0",x"00", -- 0x1568
    x"20",x"BA",x"BA",x"4C",x"20",x"B0",x"20",x"0C", -- 0x1570
    x"B0",x"A9",x"00",x"8D",x"1A",x"1C",x"8D",x"06", -- 0x1578
    x"1C",x"8D",x"04",x"1C",x"8D",x"03",x"1C",x"8D", -- 0x1580
    x"01",x"1C",x"8D",x"15",x"1C",x"8D",x"08",x"1C", -- 0x1588
    x"A9",x"02",x"20",x"3A",x"B0",x"38",x"E9",x"01", -- 0x1590
    x"A2",x"83",x"20",x"63",x"B0",x"18",x"69",x"13", -- 0x1598
    x"8D",x"00",x"1C",x"A9",x"02",x"20",x"3A",x"B0", -- 0x15A0
    x"38",x"E9",x"01",x"A2",x"20",x"20",x"63",x"B0", -- 0x15A8
    x"18",x"69",x"70",x"8D",x"02",x"1C",x"A9",x"28", -- 0x15B0
    x"8D",x"07",x"1C",x"8D",x"05",x"1C",x"AD",x"00", -- 0x15B8
    x"1C",x"18",x"E9",x"58",x"B0",x"04",x"A9",x"00", -- 0x15C0
    x"F0",x"02",x"A9",x"FF",x"D0",x"03",x"4C",x"D6", -- 0x15C8
    x"B5",x"A0",x"00",x"20",x"6E",x"BF",x"A0",x"00", -- 0x15D0
    x"20",x"26",x"BC",x"A0",x"00",x"20",x"FB",x"BB", -- 0x15D8
    x"A9",x"03",x"20",x"3A",x"B0",x"8D",x"1B",x"1C", -- 0x15E0
    x"AD",x"3B",x"1C",x"38",x"ED",x"1B",x"1C",x"8D", -- 0x15E8
    x"09",x"1C",x"AD",x"25",x"1C",x"8D",x"19",x"1C", -- 0x15F0
    x"AD",x"22",x"1C",x"8D",x"18",x"1C",x"AD",x"0C", -- 0x15F8
    x"1C",x"A8",x"B9",x"3E",x"1C",x"2D",x"0F",x"1C", -- 0x1600
    x"2D",x"12",x"1C",x"D0",x"03",x"4C",x"1B",x"B6", -- 0x1608
    x"A9",x"09",x"A0",x"02",x"91",x"01",x"A0",x"00", -- 0x1610
    x"20",x"BA",x"BA",x"A9",x"0B",x"A0",x"02",x"91", -- 0x1618
    x"01",x"AD",x"12",x"1C",x"49",x"FF",x"29",x"80", -- 0x1620
    x"48",x"AD",x"0C",x"1C",x"A8",x"B9",x"3E",x"1C", -- 0x1628
    x"49",x"FF",x"29",x"40",x"85",x"60",x"68",x"05", -- 0x1630
    x"60",x"0D",x"0C",x"1C",x"A0",x"03",x"91",x"01", -- 0x1638
    x"AD",x"00",x"1C",x"C8",x"91",x"01",x"AD",x"02", -- 0x1640
    x"1C",x"C8",x"91",x"01",x"A0",x"00",x"20",x"BA", -- 0x1648
    x"BA",x"AD",x"0C",x"1C",x"48",x"A9",x"FF",x"AA", -- 0x1650
    x"68",x"A8",x"8A",x"99",x"3E",x"1C",x"4C",x"20", -- 0x1658
    x"B0",x"20",x"0C",x"B0",x"AD",x"01",x"1C",x"18", -- 0x1660
    x"6D",x"05",x"1C",x"8D",x"01",x"1C",x"AD",x"00", -- 0x1668
    x"1C",x"6D",x"04",x"1C",x"8D",x"00",x"1C",x"AD", -- 0x1670
    x"04",x"1C",x"C9",x"80",x"90",x"04",x"A9",x"00", -- 0x1678
    x"F0",x"02",x"A9",x"FF",x"8D",x"0A",x"1C",x"AD", -- 0x1680
    x"03",x"1C",x"18",x"6D",x"07",x"1C",x"8D",x"03", -- 0x1688
    x"1C",x"AD",x"02",x"1C",x"6D",x"06",x"1C",x"8D", -- 0x1690
    x"02",x"1C",x"AD",x"06",x"1C",x"C9",x"80",x"90", -- 0x1698
    x"04",x"A9",x"00",x"F0",x"02",x"A9",x"FF",x"8D", -- 0x16A0
    x"0B",x"1C",x"AD",x"07",x"1C",x"18",x"6D",x"19", -- 0x16A8
    x"1C",x"8D",x"07",x"1C",x"AD",x"06",x"1C",x"6D", -- 0x16B0
    x"18",x"1C",x"8D",x"06",x"1C",x"AD",x"02",x"1C", -- 0x16B8
    x"18",x"E9",x"B0",x"B0",x"04",x"A9",x"00",x"F0", -- 0x16C0
    x"02",x"A9",x"FF",x"2D",x"0B",x"1C",x"D0",x"03", -- 0x16C8
    x"4C",x"61",x"B8",x"AD",x"0D",x"1C",x"D0",x"03", -- 0x16D0
    x"4C",x"ED",x"B6",x"AD",x"00",x"1C",x"38",x"ED", -- 0x16D8
    x"0E",x"1C",x"18",x"69",x"04",x"4A",x"4A",x"8D", -- 0x16E0
    x"13",x"1C",x"4C",x"05",x"B7",x"A9",x"03",x"48", -- 0x16E8
    x"AD",x"00",x"1C",x"38",x"ED",x"0E",x"1C",x"38", -- 0x16F0
    x"E9",x"0E",x"4A",x"4A",x"38",x"85",x"60",x"68", -- 0x16F8
    x"E5",x"60",x"8D",x"13",x"1C",x"AD",x"13",x"1C", -- 0x1700
    x"C9",x"04",x"90",x"04",x"A9",x"00",x"F0",x"02", -- 0x1708
    x"A9",x"FF",x"D0",x"03",x"4C",x"49",x"B8",x"AD", -- 0x1710
    x"13",x"1C",x"A8",x"B9",x"2C",x"1C",x"48",x"A9", -- 0x1718
    x"1E",x"20",x"3A",x"B0",x"18",x"85",x"60",x"68", -- 0x1720
    x"65",x"60",x"8D",x"05",x"1C",x"AD",x"13",x"1C", -- 0x1728
    x"A8",x"B9",x"28",x"1C",x"8D",x"04",x"1C",x"AD", -- 0x1730
    x"13",x"1C",x"A8",x"B9",x"34",x"1C",x"48",x"AD", -- 0x1738
    x"08",x"1C",x"A8",x"B9",x"3B",x"1C",x"38",x"ED", -- 0x1740
    x"09",x"1C",x"18",x"6D",x"1A",x"1C",x"38",x"ED", -- 0x1748
    x"1B",x"1C",x"48",x"A9",x"14",x"20",x"3A",x"B0", -- 0x1750
    x"18",x"69",x"14",x"AA",x"68",x"20",x"63",x"B0", -- 0x1758
    x"18",x"85",x"60",x"68",x"65",x"60",x"8D",x"07", -- 0x1760
    x"1C",x"AD",x"13",x"1C",x"A8",x"B9",x"30",x"1C", -- 0x1768
    x"48",x"A5",x"5E",x"29",x"01",x"85",x"60",x"68", -- 0x1770
    x"65",x"60",x"8D",x"06",x"1C",x"A0",x"00",x"20", -- 0x1778
    x"D4",x"BF",x"A9",x"02",x"38",x"ED",x"08",x"1C", -- 0x1780
    x"D0",x"03",x"4C",x"CB",x"B7",x"A9",x"01",x"8D", -- 0x1788
    x"16",x"1C",x"A9",x"02",x"38",x"ED",x"08",x"1C", -- 0x1790
    x"48",x"AD",x"04",x"1C",x"AA",x"0A",x"8A",x"6A", -- 0x1798
    x"8D",x"04",x"1C",x"AD",x"05",x"1C",x"6A",x"8D", -- 0x17A0
    x"05",x"1C",x"AD",x"06",x"1C",x"4A",x"09",x"80", -- 0x17A8
    x"8D",x"06",x"1C",x"AD",x"07",x"1C",x"6A",x"8D", -- 0x17B0
    x"07",x"1C",x"BA",x"E8",x"AD",x"16",x"1C",x"DD", -- 0x17B8
    x"00",x"01",x"B0",x"06",x"EE",x"16",x"1C",x"4C", -- 0x17C0
    x"99",x"B7",x"9A",x"AD",x"06",x"1C",x"C9",x"FA", -- 0x17C8
    x"90",x"04",x"A9",x"00",x"F0",x"02",x"A9",x"FF", -- 0x17D0
    x"D0",x"03",x"4C",x"E2",x"B7",x"A9",x"FA",x"8D", -- 0x17D8
    x"06",x"1C",x"AD",x"0E",x"1C",x"48",x"AD",x"0D", -- 0x17E0
    x"1C",x"29",x"01",x"A2",x"18",x"20",x"63",x"B0", -- 0x17E8
    x"18",x"85",x"60",x"68",x"65",x"60",x"8D",x"00", -- 0x17F0
    x"1C",x"AD",x"0D",x"1C",x"D0",x"03",x"4C",x"06", -- 0x17F8
    x"B8",x"A0",x"00",x"20",x"8B",x"BF",x"A9",x"B0", -- 0x1800
    x"8D",x"02",x"1C",x"AD",x"0D",x"1C",x"49",x"FF", -- 0x1808
    x"8D",x"0D",x"1C",x"A9",x"01",x"A0",x"02",x"91", -- 0x1810
    x"01",x"A0",x"00",x"20",x"23",x"BF",x"AD",x"1A", -- 0x1818
    x"1C",x"18",x"69",x"01",x"8D",x"1A",x"1C",x"AD", -- 0x1820
    x"08",x"1C",x"A8",x"B9",x"25",x"1C",x"8D",x"19", -- 0x1828
    x"1C",x"AD",x"08",x"1C",x"A8",x"B9",x"22",x"1C", -- 0x1830
    x"8D",x"18",x"1C",x"A9",x"0E",x"A0",x"02",x"91", -- 0x1838
    x"01",x"A0",x"00",x"20",x"BA",x"BA",x"4C",x"61", -- 0x1840
    x"B8",x"AD",x"02",x"1C",x"18",x"E9",x"B8",x"B0", -- 0x1848
    x"04",x"A9",x"00",x"F0",x"02",x"A9",x"FF",x"D0", -- 0x1850
    x"03",x"4C",x"61",x"B8",x"A9",x"FF",x"8D",x"15", -- 0x1858
    x"1C",x"AD",x"15",x"1C",x"49",x"FF",x"D0",x"03", -- 0x1860
    x"4C",x"9C",x"B8",x"A9",x"00",x"A0",x"02",x"91", -- 0x1868
    x"01",x"AD",x"0B",x"1C",x"48",x"AD",x"02",x"1C", -- 0x1870
    x"18",x"E9",x"96",x"B0",x"04",x"A9",x"00",x"F0", -- 0x1878
    x"02",x"A9",x"FF",x"85",x"60",x"68",x"25",x"60", -- 0x1880
    x"C8",x"91",x"01",x"AD",x"00",x"1C",x"C8",x"91", -- 0x1888
    x"01",x"AD",x"02",x"1C",x"C8",x"91",x"01",x"A0", -- 0x1890
    x"00",x"20",x"BA",x"BA",x"A9",x"00",x"A0",x"02", -- 0x1898
    x"91",x"01",x"A0",x"00",x"20",x"0C",x"BF",x"8D", -- 0x18A0
    x"14",x"1C",x"A9",x"FF",x"48",x"AD",x"14",x"1C", -- 0x18A8
    x"C9",x"50",x"F0",x"04",x"A9",x"00",x"F0",x"02", -- 0x18B0
    x"A9",x"FF",x"48",x"AD",x"0A",x"1C",x"49",x"FF", -- 0x18B8
    x"85",x"60",x"68",x"25",x"60",x"85",x"60",x"68", -- 0x18C0
    x"C5",x"60",x"F0",x"03",x"4C",x"D7",x"B8",x"A0", -- 0x18C8
    x"00",x"20",x"59",x"BF",x"4C",x"B7",x"BA",x"48", -- 0x18D0
    x"AD",x"14",x"1C",x"C9",x"51",x"F0",x"04",x"A9", -- 0x18D8
    x"00",x"F0",x"02",x"A9",x"FF",x"2D",x"0A",x"1C", -- 0x18E0
    x"85",x"60",x"68",x"C5",x"60",x"F0",x"03",x"4C", -- 0x18E8
    x"FA",x"B8",x"A0",x"00",x"20",x"6E",x"BF",x"4C", -- 0x18F0
    x"B7",x"BA",x"48",x"AD",x"14",x"1C",x"C9",x"52", -- 0x18F8
    x"F0",x"04",x"A9",x"00",x"F0",x"02",x"A9",x"FF", -- 0x1900
    x"48",x"AD",x"0B",x"1C",x"49",x"FF",x"85",x"60", -- 0x1908
    x"68",x"25",x"60",x"85",x"60",x"68",x"C5",x"60", -- 0x1910
    x"F0",x"03",x"4C",x"25",x"B9",x"A0",x"00",x"20", -- 0x1918
    x"A2",x"BF",x"4C",x"B7",x"BA",x"48",x"AD",x"14", -- 0x1920
    x"1C",x"C9",x"5B",x"F0",x"04",x"A9",x"00",x"F0", -- 0x1928
    x"02",x"A9",x"FF",x"2D",x"0B",x"1C",x"85",x"60", -- 0x1930
    x"68",x"C5",x"60",x"F0",x"03",x"4C",x"53",x"B9", -- 0x1938
    x"A9",x"FF",x"8D",x"06",x"1C",x"A9",x"32",x"20", -- 0x1940
    x"3A",x"B0",x"18",x"69",x"64",x"8D",x"07",x"1C", -- 0x1948
    x"4C",x"B7",x"BA",x"48",x"AD",x"14",x"1C",x"C9", -- 0x1950
    x"60",x"F0",x"04",x"A9",x"00",x"F0",x"02",x"A9", -- 0x1958
    x"FF",x"85",x"60",x"68",x"C5",x"60",x"F0",x"03", -- 0x1960
    x"4C",x"B7",x"BA",x"A9",x"02",x"A0",x"02",x"91", -- 0x1968
    x"01",x"A0",x"00",x"20",x"0C",x"BF",x"8D",x"13", -- 0x1970
    x"1C",x"AD",x"1A",x"1C",x"D0",x"03",x"4C",x"CA", -- 0x1978
    x"B9",x"AD",x"09",x"1C",x"8D",x"16",x"1C",x"AD", -- 0x1980
    x"09",x"1C",x"38",x"ED",x"13",x"1C",x"8D",x"09", -- 0x1988
    x"1C",x"AD",x"09",x"1C",x"18",x"ED",x"16",x"1C", -- 0x1990
    x"B0",x"04",x"A9",x"00",x"F0",x"02",x"A9",x"FF", -- 0x1998
    x"D0",x"03",x"4C",x"CA",x"B9",x"AD",x"08",x"1C", -- 0x19A0
    x"A8",x"B9",x"38",x"1C",x"8D",x"08",x"1C",x"A9", -- 0x19A8
    x"03",x"20",x"3A",x"B0",x"8D",x"1B",x"1C",x"AD", -- 0x19B0
    x"08",x"1C",x"A8",x"B9",x"3B",x"1C",x"38",x"ED", -- 0x19B8
    x"1B",x"1C",x"8D",x"09",x"1C",x"A9",x"00",x"8D", -- 0x19C0
    x"1A",x"1C",x"AD",x"13",x"1C",x"29",x"01",x"D0", -- 0x19C8
    x"03",x"4C",x"DE",x"B9",x"A0",x"00",x"20",x"8B", -- 0x19D0
    x"BF",x"A0",x"00",x"20",x"D4",x"BF",x"AD",x"05", -- 0x19D8
    x"1C",x"48",x"A9",x"3D",x"20",x"3A",x"B0",x"18", -- 0x19E0
    x"85",x"60",x"68",x"65",x"60",x"8D",x"05",x"1C", -- 0x19E8
    x"AD",x"04",x"1C",x"69",x"00",x"8D",x"04",x"1C", -- 0x19F0
    x"AD",x"05",x"1C",x"38",x"E9",x"1F",x"8D",x"05", -- 0x19F8
    x"1C",x"AD",x"04",x"1C",x"E9",x"00",x"8D",x"04", -- 0x1A00
    x"1C",x"A9",x"00",x"8D",x"13",x"1C",x"A9",x"02", -- 0x1A08
    x"48",x"AD",x"13",x"1C",x"18",x"69",x"03",x"A0", -- 0x1A10
    x"02",x"91",x"01",x"A0",x"00",x"20",x"0C",x"BF", -- 0x1A18
    x"2D",x"12",x"1C",x"D0",x"03",x"4C",x"8F",x"BA", -- 0x1A20
    x"AD",x"13",x"1C",x"C9",x"00",x"F0",x"04",x"A9", -- 0x1A28
    x"00",x"F0",x"02",x"A9",x"FF",x"48",x"AD",x"0C", -- 0x1A30
    x"1C",x"A8",x"B9",x"3E",x"1C",x"85",x"60",x"68", -- 0x1A38
    x"25",x"60",x"D0",x"03",x"4C",x"5F",x"BA",x"A9", -- 0x1A40
    x"15",x"A0",x"02",x"91",x"01",x"A0",x"00",x"20", -- 0x1A48
    x"BA",x"BA",x"AD",x"0C",x"1C",x"48",x"A9",x"00", -- 0x1A50
    x"AA",x"68",x"A8",x"8A",x"99",x"3E",x"1C",x"A9", -- 0x1A58
    x"14",x"A0",x"02",x"91",x"01",x"AD",x"13",x"1C", -- 0x1A60
    x"C8",x"91",x"01",x"A0",x"00",x"20",x"BA",x"BA", -- 0x1A68
    x"AD",x"0B",x"1C",x"49",x"FF",x"D0",x"03",x"4C", -- 0x1A70
    x"7F",x"BA",x"A9",x"00",x"8D",x"06",x"1C",x"AD", -- 0x1A78
    x"13",x"1C",x"A8",x"B9",x"40",x"1C",x"A0",x"02", -- 0x1A80
    x"91",x"01",x"A0",x"00",x"20",x"23",x"BF",x"BA", -- 0x1A88
    x"E8",x"AD",x"13",x"1C",x"DD",x"00",x"01",x"B0", -- 0x1A90
    x"06",x"EE",x"13",x"1C",x"4C",x"11",x"BA",x"9A", -- 0x1A98
    x"A9",x"01",x"A0",x"04",x"91",x"01",x"A0",x"02", -- 0x1AA0
    x"20",x"0C",x"BF",x"A0",x"02",x"91",x"01",x"A0", -- 0x1AA8
    x"00",x"20",x"23",x"BF",x"4C",x"B7",x"BA",x"4C", -- 0x1AB0
    x"20",x"B0",x"20",x"0C",x"B0",x"A9",x"A0",x"48", -- 0x1AB8
    x"A9",x"10",x"48",x"A0",x"00",x"B1",x"01",x"0A", -- 0x1AC0
    x"18",x"85",x"60",x"68",x"65",x"60",x"18",x"69", -- 0x1AC8
    x"01",x"85",x"34",x"68",x"85",x"35",x"B1",x"34", -- 0x1AD0
    x"A0",x"06",x"91",x"01",x"A9",x"A0",x"48",x"A9", -- 0x1AD8
    x"10",x"48",x"A0",x"00",x"B1",x"01",x"0A",x"18", -- 0x1AE0
    x"85",x"60",x"68",x"65",x"60",x"85",x"34",x"68", -- 0x1AE8
    x"85",x"35",x"B1",x"34",x"A0",x"07",x"91",x"01", -- 0x1AF0
    x"A0",x"01",x"B1",x"01",x"A0",x"08",x"91",x"01", -- 0x1AF8
    x"A0",x"02",x"B1",x"01",x"A0",x"09",x"91",x"01", -- 0x1B00
    x"A0",x"03",x"B1",x"01",x"A0",x"0A",x"91",x"01", -- 0x1B08
    x"A0",x"04",x"20",x"5E",x"B1",x"4C",x"20",x"B0", -- 0x1B10
    x"20",x"0C",x"B0",x"A0",x"00",x"20",x"FB",x"BB", -- 0x1B18
    x"A9",x"0D",x"A0",x"02",x"91",x"01",x"A0",x"00", -- 0x1B20
    x"20",x"BA",x"BA",x"A0",x"00",x"20",x"61",x"B6", -- 0x1B28
    x"A9",x"11",x"A0",x"02",x"91",x"01",x"A0",x"00", -- 0x1B30
    x"20",x"BA",x"BA",x"A9",x"05",x"A0",x"02",x"91", -- 0x1B38
    x"01",x"A0",x"00",x"20",x"BA",x"BA",x"AD",x"15", -- 0x1B40
    x"1C",x"F0",x"D0",x"A9",x"03",x"A0",x"02",x"91", -- 0x1B48
    x"01",x"A9",x"0F",x"C8",x"91",x"01",x"A0",x"00", -- 0x1B50
    x"20",x"2D",x"B3",x"A9",x"16",x"A0",x"02",x"91", -- 0x1B58
    x"01",x"AD",x"11",x"1C",x"C8",x"91",x"01",x"AD", -- 0x1B60
    x"10",x"1C",x"C8",x"91",x"01",x"AD",x"00",x"1C", -- 0x1B68
    x"C8",x"91",x"01",x"A0",x"00",x"20",x"BA",x"BA", -- 0x1B70
    x"AD",x"0C",x"1C",x"A8",x"B9",x"3E",x"1C",x"D0", -- 0x1B78
    x"03",x"4C",x"F8",x"BB",x"AD",x"0C",x"1C",x"48", -- 0x1B80
    x"AD",x"0C",x"1C",x"A8",x"B9",x"20",x"1C",x"38", -- 0x1B88
    x"E9",x"01",x"AA",x"68",x"A8",x"8A",x"99",x"20", -- 0x1B90
    x"1C",x"A0",x"00",x"20",x"26",x"BC",x"AD",x"0F", -- 0x1B98
    x"1C",x"2D",x"21",x"1C",x"D0",x"03",x"4C",x"F8", -- 0x1BA0
    x"BB",x"AD",x"20",x"1C",x"C9",x"00",x"F0",x"04", -- 0x1BA8
    x"A9",x"00",x"F0",x"02",x"A9",x"FF",x"D0",x"03", -- 0x1BB0
    x"4C",x"F0",x"BB",x"A9",x"02",x"A0",x"02",x"91", -- 0x1BB8
    x"01",x"A9",x"10",x"C8",x"91",x"01",x"A0",x"00", -- 0x1BC0
    x"20",x"2D",x"B3",x"A9",x"01",x"85",x"38",x"20", -- 0x1BC8
    x"F5",x"B0",x"47",x"41",x"4D",x"45",x"20",x"4F", -- 0x1BD0
    x"56",x"45",x"52",x"20",x"50",x"4C",x"41",x"59", -- 0x1BD8
    x"45",x"52",x"20",x"31",x"00",x"A9",x"FF",x"A0", -- 0x1BE0
    x"02",x"91",x"01",x"A0",x"00",x"20",x"5B",x"BE", -- 0x1BE8
    x"AD",x"0C",x"1C",x"49",x"01",x"8D",x"0C",x"1C", -- 0x1BF0
    x"4C",x"20",x"B0",x"20",x"0C",x"B0",x"A9",x"03", -- 0x1BF8
    x"A0",x"02",x"91",x"01",x"AD",x"0C",x"1C",x"C8", -- 0x1C00
    x"91",x"01",x"AD",x"0D",x"1C",x"C8",x"91",x"01", -- 0x1C08
    x"A0",x"00",x"20",x"BA",x"BA",x"A9",x"00",x"A0", -- 0x1C10
    x"02",x"91",x"01",x"A0",x"00",x"20",x"0C",x"BF", -- 0x1C18
    x"8D",x"0E",x"1C",x"4C",x"20",x"B0",x"20",x"0C", -- 0x1C20
    x"B0",x"AD",x"12",x"1C",x"D0",x"03",x"4C",x"69", -- 0x1C28
    x"BC",x"A9",x"07",x"A0",x"02",x"91",x"01",x"AD", -- 0x1C30
    x"0C",x"1C",x"A8",x"B9",x"1E",x"1C",x"A0",x"03", -- 0x1C38
    x"91",x"01",x"AD",x"0C",x"1C",x"A8",x"B9",x"1C", -- 0x1C40
    x"1C",x"A0",x"04",x"91",x"01",x"AD",x"0C",x"1C", -- 0x1C48
    x"6A",x"6A",x"48",x"AD",x"0C",x"1C",x"A8",x"B9", -- 0x1C50
    x"20",x"1C",x"18",x"85",x"60",x"68",x"65",x"60", -- 0x1C58
    x"A0",x"05",x"91",x"01",x"A0",x"00",x"20",x"BA", -- 0x1C60
    x"BA",x"4C",x"20",x"B0",x"20",x"0C",x"B0",x"A9", -- 0x1C68
    x"00",x"8D",x"0F",x"1C",x"8D",x"12",x"1C",x"A9", -- 0x1C70
    x"19",x"A0",x"02",x"91",x"01",x"A0",x"00",x"20", -- 0x1C78
    x"BA",x"BA",x"A9",x"01",x"8D",x"13",x"1C",x"A9", -- 0x1C80
    x"90",x"48",x"A9",x"00",x"18",x"69",x"08",x"A0", -- 0x1C88
    x"00",x"85",x"34",x"68",x"85",x"35",x"B1",x"34", -- 0x1C90
    x"20",x"3A",x"B0",x"48",x"A9",x"FF",x"20",x"3A", -- 0x1C98
    x"B0",x"8D",x"16",x"1C",x"BA",x"E8",x"AD",x"13", -- 0x1CA0
    x"1C",x"DD",x"00",x"01",x"B0",x"06",x"EE",x"13", -- 0x1CA8
    x"1C",x"4C",x"9C",x"BC",x"9A",x"A9",x"0C",x"A0", -- 0x1CB0
    x"02",x"91",x"01",x"A0",x"00",x"20",x"BA",x"BA", -- 0x1CB8
    x"A9",x"00",x"A0",x"02",x"91",x"01",x"A0",x"00", -- 0x1CC0
    x"20",x"0C",x"BF",x"D0",x"03",x"4C",x"D3",x"BC", -- 0x1CC8
    x"4C",x"20",x"B0",x"A0",x"00",x"20",x"E6",x"B4", -- 0x1CD0
    x"A9",x"03",x"A0",x"02",x"91",x"01",x"A9",x"0F", -- 0x1CD8
    x"C8",x"91",x"01",x"A0",x"00",x"20",x"2D",x"B3", -- 0x1CE0
    x"A9",x"17",x"A0",x"02",x"91",x"01",x"AD",x"11", -- 0x1CE8
    x"1C",x"C8",x"91",x"01",x"AD",x"10",x"1C",x"C8", -- 0x1CF0
    x"91",x"01",x"A0",x"00",x"20",x"BA",x"BA",x"A9", -- 0x1CF8
    x"01",x"85",x"38",x"20",x"18",x"B1",x"20",x"F5", -- 0x1D00
    x"B0",x"11",x"11",x"1D",x"20",x"50",x"55",x"53", -- 0x1D08
    x"48",x"20",x"27",x"46",x"31",x"27",x"20",x"54", -- 0x1D10
    x"4F",x"20",x"42",x"45",x"47",x"49",x"4E",x"00", -- 0x1D18
    x"A9",x"1A",x"A0",x"02",x"91",x"01",x"AD",x"0E", -- 0x1D20
    x"1C",x"C8",x"91",x"01",x"AD",x"0D",x"1C",x"C8", -- 0x1D28
    x"91",x"01",x"A0",x"00",x"20",x"BA",x"BA",x"A0", -- 0x1D30
    x"00",x"20",x"76",x"B5",x"A9",x"0D",x"A0",x"02", -- 0x1D38
    x"91",x"01",x"A0",x"00",x"20",x"BA",x"BA",x"AD", -- 0x1D40
    x"0E",x"1C",x"C9",x"08",x"90",x"04",x"A9",x"00", -- 0x1D48
    x"F0",x"02",x"A9",x"FF",x"D0",x"03",x"4C",x"5E", -- 0x1D50
    x"BD",x"A9",x"08",x"8D",x"0E",x"1C",x"AD",x"0D", -- 0x1D58
    x"1C",x"D0",x"03",x"4C",x"73",x"BD",x"AD",x"00", -- 0x1D60
    x"1C",x"38",x"ED",x"0E",x"1C",x"8D",x"16",x"1C", -- 0x1D68
    x"4C",x"80",x"BD",x"AD",x"00",x"1C",x"38",x"ED", -- 0x1D70
    x"0E",x"1C",x"38",x"E9",x"17",x"8D",x"16",x"1C", -- 0x1D78
    x"A9",x"FF",x"48",x"AD",x"16",x"1C",x"C9",x"00", -- 0x1D80
    x"F0",x"04",x"A9",x"00",x"F0",x"02",x"A9",x"FF", -- 0x1D88
    x"85",x"60",x"68",x"C5",x"60",x"F0",x"03",x"4C", -- 0x1D90
    x"9D",x"BD",x"4C",x"D4",x"BD",x"48",x"AD",x"16", -- 0x1D98
    x"1C",x"C9",x"80",x"90",x"04",x"A9",x"00",x"F0", -- 0x1DA0
    x"02",x"A9",x"FF",x"85",x"60",x"68",x"C5",x"60", -- 0x1DA8
    x"F0",x"03",x"4C",x"C4",x"BD",x"A9",x"03",x"20", -- 0x1DB0
    x"3A",x"B0",x"4A",x"6D",x"0E",x"1C",x"8D",x"0E", -- 0x1DB8
    x"1C",x"4C",x"D4",x"BD",x"A9",x"03",x"20",x"3A", -- 0x1DC0
    x"B0",x"49",x"FF",x"4A",x"09",x"80",x"6D",x"0E", -- 0x1DC8
    x"1C",x"8D",x"0E",x"1C",x"A9",x"1A",x"A0",x"02", -- 0x1DD0
    x"91",x"01",x"AD",x"0E",x"1C",x"C8",x"91",x"01", -- 0x1DD8
    x"AD",x"0D",x"1C",x"C8",x"91",x"01",x"A0",x"00", -- 0x1DE0
    x"20",x"BA",x"BA",x"A0",x"00",x"20",x"61",x"B6", -- 0x1DE8
    x"A9",x"1C",x"A0",x"02",x"91",x"01",x"A0",x"00", -- 0x1DF0
    x"20",x"BA",x"BA",x"A9",x"08",x"A0",x"02",x"91", -- 0x1DF8
    x"01",x"A0",x"00",x"20",x"BA",x"BA",x"A9",x"00", -- 0x1E00
    x"A0",x"02",x"91",x"01",x"A0",x"00",x"20",x"0C", -- 0x1E08
    x"BF",x"C9",x"01",x"F0",x"04",x"A9",x"00",x"F0", -- 0x1E10
    x"02",x"A9",x"FF",x"D0",x"03",x"4C",x"23",x"BE", -- 0x1E18
    x"4C",x"20",x"B0",x"A9",x"05",x"A0",x"02",x"91", -- 0x1E20
    x"01",x"A0",x"00",x"20",x"BA",x"BA",x"AD",x"15", -- 0x1E28
    x"1C",x"D0",x"03",x"4C",x"3C",x"BD",x"A9",x"16", -- 0x1E30
    x"A0",x"02",x"91",x"01",x"A9",x"00",x"C8",x"91", -- 0x1E38
    x"01",x"A9",x"00",x"C8",x"91",x"01",x"AD",x"00", -- 0x1E40
    x"1C",x"C8",x"91",x"01",x"A0",x"00",x"20",x"BA", -- 0x1E48
    x"BA",x"A9",x"00",x"D0",x"03",x"4C",x"B5",x"BC", -- 0x1E50
    x"4C",x"20",x"B0",x"20",x"0C",x"B0",x"A9",x"01", -- 0x1E58
    x"8D",x"16",x"1C",x"A0",x"00",x"B1",x"01",x"48", -- 0x1E60
    x"A9",x"05",x"A0",x"03",x"91",x"01",x"A0",x"01", -- 0x1E68
    x"20",x"BA",x"BA",x"BA",x"E8",x"AD",x"16",x"1C", -- 0x1E70
    x"DD",x"00",x"01",x"B0",x"06",x"EE",x"16",x"1C", -- 0x1E78
    x"4C",x"68",x"BE",x"9A",x"4C",x"20",x"B0",x"20", -- 0x1E80
    x"0C",x"B0",x"A9",x"07",x"A0",x"02",x"91",x"01", -- 0x1E88
    x"A0",x"00",x"20",x"3E",x"B3",x"A9",x"01",x"85", -- 0x1E90
    x"38",x"20",x"F5",x"B0",x"93",x"11",x"11",x"2A", -- 0x1E98
    x"20",x"4E",x"55",x"4D",x"42",x"45",x"52",x"20", -- 0x1EA0
    x"4F",x"46",x"20",x"50",x"4C",x"41",x"59",x"45", -- 0x1EA8
    x"52",x"53",x"00",x"20",x"18",x"B1",x"20",x"F5", -- 0x1EB0
    x"B0",x"11",x"1D",x"1D",x"27",x"46",x"31",x"27", -- 0x1EB8
    x"20",x"2D",x"20",x"31",x"20",x"50",x"4C",x"41", -- 0x1EC0
    x"59",x"45",x"52",x"00",x"20",x"18",x"B1",x"20", -- 0x1EC8
    x"F5",x"B0",x"11",x"1D",x"1D",x"27",x"46",x"33", -- 0x1ED0
    x"27",x"20",x"2D",x"20",x"32",x"20",x"50",x"4C", -- 0x1ED8
    x"41",x"59",x"45",x"52",x"53",x"00",x"A9",x"1B", -- 0x1EE0
    x"A0",x"02",x"91",x"01",x"A0",x"00",x"20",x"BA", -- 0x1EE8
    x"BA",x"A9",x"00",x"A0",x"02",x"91",x"01",x"A0", -- 0x1EF0
    x"00",x"20",x"0C",x"BF",x"C9",x"03",x"F0",x"04", -- 0x1EF8
    x"A9",x"00",x"F0",x"02",x"A9",x"FF",x"8D",x"0F", -- 0x1F00
    x"1C",x"4C",x"20",x"B0",x"20",x"0C",x"B0",x"A9", -- 0x1F08
    x"00",x"48",x"A9",x"68",x"18",x"A0",x"00",x"71", -- 0x1F10
    x"01",x"85",x"34",x"68",x"85",x"35",x"B1",x"34", -- 0x1F18
    x"4C",x"20",x"B0",x"20",x"0C",x"B0",x"AD",x"0C", -- 0x1F20
    x"1C",x"48",x"AD",x"0C",x"1C",x"A8",x"B9",x"1E", -- 0x1F28
    x"1C",x"18",x"A0",x"00",x"71",x"01",x"AA",x"68", -- 0x1F30
    x"A8",x"8A",x"99",x"1E",x"1C",x"AD",x"0C",x"1C", -- 0x1F38
    x"48",x"AD",x"0C",x"1C",x"A8",x"B9",x"1C",x"1C", -- 0x1F40
    x"69",x"00",x"AA",x"68",x"A8",x"8A",x"99",x"1C", -- 0x1F48
    x"1C",x"A0",x"01",x"20",x"26",x"BC",x"4C",x"20", -- 0x1F50
    x"B0",x"20",x"0C",x"B0",x"AD",x"04",x"1C",x"29", -- 0x1F58
    x"80",x"D0",x"03",x"4C",x"6B",x"BF",x"A0",x"00", -- 0x1F60
    x"20",x"8B",x"BF",x"4C",x"20",x"B0",x"20",x"0C", -- 0x1F68
    x"B0",x"AD",x"04",x"1C",x"C9",x"80",x"90",x"04", -- 0x1F70
    x"A9",x"00",x"F0",x"02",x"A9",x"FF",x"D0",x"03", -- 0x1F78
    x"4C",x"88",x"BF",x"A0",x"00",x"20",x"8B",x"BF", -- 0x1F80
    x"4C",x"20",x"B0",x"20",x"0C",x"B0",x"A9",x"00", -- 0x1F88
    x"38",x"ED",x"05",x"1C",x"8D",x"05",x"1C",x"A9", -- 0x1F90
    x"00",x"ED",x"04",x"1C",x"8D",x"04",x"1C",x"4C", -- 0x1F98
    x"20",x"B0",x"20",x"0C",x"B0",x"AD",x"06",x"1C", -- 0x1FA0
    x"29",x"80",x"D0",x"03",x"4C",x"B4",x"BF",x"A0", -- 0x1FA8
    x"00",x"20",x"D4",x"BF",x"4C",x"20",x"B0",x"20", -- 0x1FB0
    x"0C",x"B0",x"AD",x"06",x"1C",x"C9",x"80",x"90", -- 0x1FB8
    x"04",x"A9",x"00",x"F0",x"02",x"A9",x"FF",x"D0", -- 0x1FC0
    x"03",x"4C",x"D1",x"BF",x"A0",x"00",x"20",x"D4", -- 0x1FC8
    x"BF",x"4C",x"20",x"B0",x"20",x"0C",x"B0",x"A9", -- 0x1FD0
    x"00",x"38",x"ED",x"07",x"1C",x"8D",x"07",x"1C", -- 0x1FD8
    x"A9",x"00",x"ED",x"06",x"1C",x"8D",x"06",x"1C", -- 0x1FE0
    x"4C",x"20",x"B0",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x1FE8
    x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x1FF0
    x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"00"  -- 0x1FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
