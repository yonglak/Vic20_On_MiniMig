-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity cart_rom is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of cart_rom is


  type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"F2",x"B6",x"B3",x"B2",x"41",x"30",x"C3",x"C2", -- 0x0000
	-- x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C2", -- 0x0000 -- test
    x"CD",x"A9",x"1E",x"8D",x"0F",x"90",x"A9",x"20", -- 0x0008
    x"85",x"8B",x"A9",x"00",x"20",x"7B",x"B1",x"A0", -- 0x0010
    x"0F",x"B9",x"F4",x"BB",x"99",x"B0",x"1E",x"A9", -- 0x0018
    x"02",x"99",x"B0",x"96",x"A9",x"06",x"99",x"8C", -- 0x0020
    x"97",x"99",x"B8",x"97",x"B9",x"04",x"BC",x"99", -- 0x0028
    x"DD",x"1E",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x0030
    x"B9",x"14",x"BC",x"99",x"8C",x"1F",x"B9",x"24", -- 0x0038
    x"BC",x"99",x"B8",x"1F",x"88",x"10",x"D2",x"A0", -- 0x0040
    x"2C",x"A9",x"1F",x"85",x"8A",x"A2",x"01",x"86", -- 0x0048
    x"87",x"86",x"86",x"86",x"88",x"8E",x"27",x"18", -- 0x0050
    x"CA",x"86",x"7D",x"A5",x"7D",x"F0",x"FC",x"C6", -- 0x0058
    x"7D",x"C6",x"87",x"D0",x"F6",x"A9",x"05",x"85", -- 0x0060
    x"87",x"E6",x"88",x"A5",x"88",x"4A",x"4A",x"B0", -- 0x0068
    x"17",x"A9",x"22",x"8D",x"38",x"1F",x"8D",x"3F", -- 0x0070
    x"1F",x"A2",x"05",x"BD",x"0F",x"1E",x"29",x"7F", -- 0x0078
    x"9D",x"39",x"1F",x"CA",x"10",x"F5",x"30",x"0A", -- 0x0080
    x"A9",x"20",x"A2",x"07",x"9D",x"38",x"1F",x"CA", -- 0x0088
    x"10",x"FA",x"CE",x"27",x"18",x"D0",x"13",x"A9", -- 0x0090
    x"03",x"8D",x"27",x"18",x"98",x"48",x"A4",x"8A", -- 0x0098
    x"B9",x"D1",x"BD",x"8D",x"0B",x"90",x"C6",x"8A", -- 0x00A0
    x"68",x"A8",x"C6",x"86",x"D0",x"AD",x"B9",x"77", -- 0x00A8
    x"BD",x"8D",x"0C",x"90",x"B9",x"A4",x"BD",x"85", -- 0x00B0
    x"86",x"88",x"10",x"9F",x"C8",x"8C",x"0B",x"90", -- 0x00B8
    x"4C",x"C4",x"B2",x"AD",x"0E",x"90",x"29",x"F0", -- 0x00C0
    x"8D",x"0E",x"90",x"20",x"29",x"A2",x"A2",x"0B", -- 0x00C8
    x"BD",x"B5",x"A2",x"9D",x"86",x"1E",x"CA",x"10", -- 0x00D0
    x"F7",x"A2",x"0F",x"BD",x"28",x"A3",x"9D",x"E5", -- 0x00D8
    x"1F",x"CA",x"10",x"F7",x"A9",x"28",x"85",x"28", -- 0x00E0
    x"A9",x"B0",x"85",x"EF",x"A9",x"1E",x"85",x"F0", -- 0x00E8
    x"A9",x"C6",x"85",x"F1",x"A9",x"1E",x"85",x"F2", -- 0x00F0
    x"A2",x"03",x"A9",x"36",x"85",x"20",x"BD",x"3B", -- 0x00F8
    x"A3",x"85",x"EB",x"BD",x"43",x"A3",x"85",x"EC", -- 0x0100
    x"BD",x"3F",x"A3",x"85",x"ED",x"BD",x"47",x"A3", -- 0x0108
    x"85",x"EE",x"8A",x"48",x"A9",x"13",x"8D",x"38", -- 0x0110
    x"18",x"8D",x"36",x"18",x"A5",x"7D",x"F0",x"FC", -- 0x0118
    x"C6",x"7D",x"CE",x"36",x"18",x"D0",x"F5",x"A9", -- 0x0120
    x"03",x"8D",x"36",x"18",x"20",x"5B",x"A5",x"C6", -- 0x0128
    x"20",x"AD",x"38",x"18",x"30",x"1F",x"AC",x"38", -- 0x0130
    x"18",x"C0",x"12",x"B0",x"12",x"A9",x"20",x"91", -- 0x0138
    x"EF",x"91",x"F1",x"C0",x"11",x"B0",x"08",x"B1", -- 0x0140
    x"EB",x"91",x"EF",x"B1",x"ED",x"91",x"F1",x"CE", -- 0x0148
    x"38",x"18",x"4C",x"1C",x"A1",x"A2",x"14",x"20", -- 0x0150
    x"C6",x"B2",x"A5",x"EF",x"18",x"69",x"2C",x"85", -- 0x0158
    x"EF",x"90",x"02",x"E6",x"F0",x"A5",x"F1",x"18", -- 0x0160
    x"69",x"2C",x"85",x"F1",x"90",x"02",x"E6",x"F2", -- 0x0168
    x"E6",x"28",x"E6",x"28",x"68",x"AA",x"CA",x"10", -- 0x0170
    x"81",x"20",x"C4",x"B2",x"A9",x"52",x"85",x"87", -- 0x0178
    x"A2",x"03",x"BC",x"43",x"BC",x"A5",x"87",x"99", -- 0x0180
    x"90",x"1F",x"A9",x"05",x"99",x"90",x"97",x"C6", -- 0x0188
    x"87",x"BD",x"37",x"A3",x"9D",x"96",x"1F",x"CA", -- 0x0190
    x"D0",x"E8",x"86",x"87",x"86",x"88",x"A9",x"09", -- 0x0198
    x"85",x"8B",x"20",x"D0",x"B2",x"4A",x"85",x"8B", -- 0x01A0
    x"E6",x"8B",x"A0",x"03",x"A9",x"20",x"99",x"92", -- 0x01A8
    x"1F",x"A9",x"00",x"99",x"92",x"97",x"88",x"10", -- 0x01B0
    x"F3",x"8D",x"AA",x"97",x"8D",x"AB",x"97",x"A9", -- 0x01B8
    x"20",x"8D",x"AA",x"1F",x"8D",x"AB",x"1F",x"A2", -- 0x01C0
    x"1E",x"20",x"C6",x"B2",x"A5",x"87",x"F8",x"69", -- 0x01C8
    x"01",x"85",x"87",x"D8",x"A5",x"87",x"C5",x"8B", -- 0x01D0
    x"D0",x"09",x"E6",x"88",x"A9",x"53",x"8D",x"A7", -- 0x01D8
    x"1F",x"D0",x"04",x"A9",x"20",x"D0",x"F7",x"A9", -- 0x01E0
    x"30",x"8D",x"94",x"1F",x"8D",x"95",x"1F",x"A5", -- 0x01E8
    x"87",x"29",x"0F",x"09",x"30",x"8D",x"93",x"1F", -- 0x01F0
    x"A5",x"87",x"29",x"F0",x"F0",x"05",x"A9",x"31", -- 0x01F8
    x"8D",x"92",x"1F",x"A5",x"88",x"F0",x"0A",x"A9", -- 0x0200
    x"18",x"8D",x"AA",x"1F",x"A9",x"32",x"8D",x"AB", -- 0x0208
    x"1F",x"A2",x"1E",x"20",x"C6",x"B2",x"A5",x"87", -- 0x0210
    x"C9",x"10",x"D0",x"8E",x"A2",x"78",x"20",x"C6", -- 0x0218
    x"B2",x"AD",x"43",x"18",x"D0",x"23",x"4C",x"AB", -- 0x0220
    x"A3",x"A9",x"2D",x"85",x"90",x"85",x"91",x"A9", -- 0x0228
    x"36",x"85",x"20",x"A9",x"03",x"85",x"40",x"A9", -- 0x0230
    x"00",x"85",x"7F",x"A9",x"7E",x"8D",x"0F",x"90", -- 0x0238
    x"A9",x"20",x"85",x"8B",x"58",x"EA",x"4C",x"79", -- 0x0240
    x"B1",x"A9",x"20",x"85",x"8B",x"20",x"79",x"B1", -- 0x0248
    x"A9",x"3E",x"8D",x"0F",x"90",x"20",x"C4",x"B2", -- 0x0250
    x"A9",x"4B",x"85",x"80",x"A9",x"A3",x"85",x"81", -- 0x0258
    x"A9",x"B1",x"85",x"82",x"A9",x"1E",x"85",x"83", -- 0x0260
    x"A9",x"06",x"85",x"87",x"A0",x"0F",x"B1",x"80", -- 0x0268
    x"29",x"3F",x"91",x"82",x"88",x"10",x"F7",x"20", -- 0x0270
    x"C4",x"B2",x"A5",x"80",x"18",x"69",x"10",x"85", -- 0x0278
    x"80",x"90",x"02",x"E6",x"81",x"A5",x"82",x"18", -- 0x0280
    x"69",x"2C",x"85",x"82",x"90",x"02",x"E6",x"83", -- 0x0288
    x"C6",x"87",x"D0",x"D8",x"A9",x"17",x"85",x"87", -- 0x0290
    x"A5",x"87",x"29",x"07",x"A0",x"0C",x"99",x"0B", -- 0x0298
    x"97",x"88",x"10",x"FA",x"A2",x"0C",x"20",x"C6", -- 0x02A0
    x"B2",x"C6",x"87",x"10",x"EB",x"A2",x"96",x"20", -- 0x02A8
    x"C6",x"B2",x"4C",x"AB",x"A3",x"16",x"09",x"03", -- 0x02B0
    x"20",x"12",x"01",x"14",x"20",x"12",x"01",x"03", -- 0x02B8
    x"05",x"20",x"2D",x"09",x"0E",x"13",x"14",x"12", -- 0x02C0
    x"15",x"03",x"14",x"09",x"0F",x"0E",x"13",x"2D", -- 0x02C8
    x"20",x"20",x"04",x"0F",x"04",x"07",x"05",x"20", -- 0x02D0
    x"03",x"01",x"14",x"13",x"20",x"01",x"0E",x"04", -- 0x02D8
    x"20",x"20",x"12",x"05",x"04",x"20",x"12",x"01", -- 0x02E0
    x"14",x"13",x"20",x"14",x"0F",x"20",x"05",x"01", -- 0x02E8
    x"14",x"20",x"14",x"09",x"0D",x"05",x"20",x"12", -- 0x02F0
    x"15",x"0E",x"13",x"20",x"0F",x"15",x"14",x"2E", -- 0x02F8
    x"20",x"20",x"31",x"30",x"20",x"03",x"08",x"05", -- 0x0300
    x"05",x"13",x"05",x"13",x"20",x"02",x"05",x"06", -- 0x0308
    x"0F",x"12",x"05",x"20",x"20",x"20",x"20",x"20", -- 0x0310
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x0318
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x0320
    x"10",x"15",x"13",x"08",x"20",x"86",x"B1",x"20", -- 0x0328
    x"14",x"0F",x"20",x"13",x"14",x"01",x"12",x"14", -- 0x0330
    x"10",x"14",x"13",x"13",x"13",x"D1",x"C1",x"F1", -- 0x0338
    x"02",x"E1",x"13",x"A3",x"A3",x"A2",x"A2",x"A2", -- 0x0340
    x"A3",x"A2",x"A3",x"54",x"48",x"49",x"53",x"20", -- 0x0348
    x"50",x"52",x"4F",x"47",x"52",x"41",x"4D",x"20", -- 0x0350
    x"57",x"41",x"53",x"20",x"20",x"20",x"43",x"52", -- 0x0358
    x"45",x"41",x"54",x"45",x"44",x"20",x"42",x"59", -- 0x0360
    x"20",x"20",x"20",x"20",x"2D",x"42",x"49",x"4C", -- 0x0368
    x"4C",x"20",x"48",x"49",x"4E",x"44",x"4F",x"52", -- 0x0370
    x"46",x"46",x"2D",x"20",x"20",x"20",x"4E",x"4F", -- 0x0378
    x"56",x"2E",x"20",x"35",x"2C",x"20",x"31",x"39", -- 0x0380
    x"38",x"31",x"20",x"20",x"20",x"56",x"49",x"43", -- 0x0388
    x"20",x"43",x"4F",x"4D",x"4D",x"41",x"4E",x"44", -- 0x0390
    x"4F",x"53",x"20",x"20",x"20",x"4B",x"2E",x"20", -- 0x0398
    x"4F",x"46",x"20",x"50",x"2E",x"2C",x"20",x"55", -- 0x03A0
    x"53",x"41",x"20",x"A9",x"CE",x"8D",x"0F",x"90", -- 0x03A8
    x"A2",x"06",x"86",x"7E",x"A2",x"01",x"86",x"9F", -- 0x03B0
    x"86",x"E0",x"CA",x"86",x"E1",x"20",x"CD",x"B8", -- 0x03B8
    x"20",x"00",x"B0",x"20",x"C4",x"B2",x"A9",x"12", -- 0x03C0
    x"8D",x"42",x"18",x"A9",x"00",x"85",x"E3",x"A9", -- 0x03C8
    x"02",x"8D",x"26",x"18",x"A5",x"7D",x"F0",x"FC", -- 0x03D0
    x"C6",x"9E",x"D0",x"11",x"A5",x"7E",x"85",x"9E", -- 0x03D8
    x"8D",x"41",x"18",x"20",x"69",x"AB",x"20",x"A1", -- 0x03E0
    x"B8",x"A5",x"9D",x"D0",x"25",x"AD",x"0B",x"18", -- 0x03E8
    x"30",x"10",x"CE",x"0B",x"18",x"D0",x"0B",x"A4", -- 0x03F0
    x"E1",x"B9",x"00",x"BE",x"8D",x"0B",x"18",x"20", -- 0x03F8
    x"7D",x"A4",x"20",x"EC",x"AD",x"20",x"A1",x"B8", -- 0x0400
    x"A5",x"9D",x"D0",x"06",x"A9",x"00",x"85",x"7D", -- 0x0408
    x"F0",x"C2",x"20",x"5B",x"A5",x"A9",x"00",x"8D", -- 0x0410
    x"41",x"18",x"A9",x"26",x"85",x"80",x"A9",x"1F", -- 0x0418
    x"85",x"81",x"20",x"A1",x"AC",x"20",x"C4",x"B2", -- 0x0420
    x"20",x"C4",x"B2",x"4C",x"C3",x"A0",x"A9",x"00", -- 0x0428
    x"85",x"E4",x"A2",x"02",x"B5",x"20",x"38",x"E5", -- 0x0430
    x"90",x"C9",x"08",x"B0",x"13",x"B5",x"28",x"38", -- 0x0438
    x"E5",x"91",x"C9",x"08",x"B0",x"04",x"E6",x"E4", -- 0x0440
    x"D0",x"0A",x"C9",x"F8",x"B0",x"F8",x"90",x"04", -- 0x0448
    x"C9",x"F8",x"B0",x"E9",x"CA",x"10",x"DD",x"CE", -- 0x0450
    x"42",x"18",x"D0",x"20",x"A9",x"06",x"85",x"8B", -- 0x0458
    x"20",x"D0",x"B2",x"69",x"08",x"8D",x"42",x"18", -- 0x0460
    x"A9",x"04",x"85",x"8B",x"20",x"D0",x"B2",x"4A", -- 0x0468
    x"85",x"E3",x"38",x"E5",x"8D",x"4A",x"B0",x"04", -- 0x0470
    x"A9",x"FF",x"85",x"E3",x"60",x"A0",x"1F",x"A9", -- 0x0478
    x"20",x"99",x"00",x"00",x"88",x"10",x"FA",x"20", -- 0x0480
    x"5B",x"A5",x"A0",x"1F",x"B9",x"64",x"BC",x"99", -- 0x0488
    x"00",x"00",x"88",x"10",x"F7",x"A6",x"7F",x"B5", -- 0x0490
    x"48",x"F0",x"09",x"29",x"03",x"95",x"40",x"D6", -- 0x0498
    x"48",x"4C",x"48",x"A5",x"B5",x"30",x"4A",x"90", -- 0x04A0
    x"03",x"4C",x"0E",x"A5",x"20",x"3C",x"A6",x"AD", -- 0x04A8
    x"0A",x"18",x"30",x"33",x"D5",x"38",x"F0",x"2F", -- 0x04B0
    x"B5",x"38",x"85",x"8A",x"AD",x"0A",x"18",x"95", -- 0x04B8
    x"38",x"20",x"0D",x"A6",x"08",x"A6",x"82",x"28", -- 0x04C0
    x"D0",x"19",x"A5",x"8A",x"38",x"F5",x"38",x"29", -- 0x04C8
    x"03",x"C9",x"02",x"F0",x"03",x"4C",x"41",x"A5", -- 0x04D0
    x"B5",x"38",x"E9",x"01",x"29",x"03",x"95",x"40", -- 0x04D8
    x"4C",x"45",x"A5",x"A5",x"8A",x"95",x"38",x"20", -- 0x04E0
    x"0D",x"A6",x"08",x"A6",x"82",x"28",x"F0",x"1E", -- 0x04E8
    x"F6",x"38",x"B5",x"38",x"29",x"03",x"95",x"38", -- 0x04F0
    x"20",x"0D",x"A6",x"08",x"A6",x"82",x"28",x"F0", -- 0x04F8
    x"40",x"F6",x"38",x"F6",x"38",x"B5",x"38",x"29", -- 0x0500
    x"03",x"95",x"38",x"4C",x"41",x"A5",x"B4",x"38", -- 0x0508
    x"B8",x"D0",x"04",x"D6",x"28",x"50",x"10",x"88", -- 0x0510
    x"D0",x"04",x"F6",x"20",x"50",x"09",x"88",x"D0", -- 0x0518
    x"04",x"F6",x"28",x"50",x"02",x"D6",x"20",x"F6", -- 0x0520
    x"30",x"B5",x"20",x"10",x"02",x"F6",x"20",x"C9", -- 0x0528
    x"40",x"90",x"02",x"D6",x"20",x"B5",x"28",x"10", -- 0x0530
    x"02",x"F6",x"28",x"C9",x"70",x"90",x"02",x"D6", -- 0x0538
    x"28",x"B5",x"38",x"95",x"40",x"20",x"AB",x"A6", -- 0x0540
    x"CA",x"30",x"03",x"4C",x"97",x"A4",x"AD",x"21", -- 0x0548
    x"18",x"D0",x"05",x"AD",x"22",x"18",x"D0",x"03", -- 0x0550
    x"20",x"1D",x"A7",x"A6",x"7F",x"86",x"8B",x"B5", -- 0x0558
    x"20",x"85",x"8C",x"B5",x"28",x"20",x"15",x"AB", -- 0x0560
    x"F0",x"03",x"4C",x"05",x"A6",x"B5",x"40",x"AA", -- 0x0568
    x"A5",x"82",x"F0",x"21",x"A5",x"85",x"F0",x"11", -- 0x0570
    x"B5",x"10",x"91",x"80",x"A9",x"02",x"91",x"8E", -- 0x0578
    x"A5",x"85",x"C9",x"11",x"D0",x"03",x"4C",x"05", -- 0x0580
    x"A6",x"A0",x"16",x"B5",x"14",x"91",x"80",x"A9", -- 0x0588
    x"02",x"91",x"8E",x"D0",x"70",x"A5",x"84",x"C9", -- 0x0590
    x"11",x"D0",x"1E",x"A5",x"85",x"F0",x"0E",x"B5", -- 0x0598
    x"18",x"91",x"80",x"A9",x"02",x"91",x"8E",x"A5", -- 0x05A0
    x"85",x"C9",x"11",x"F0",x"58",x"A0",x"16",x"B5", -- 0x05A8
    x"1C",x"91",x"80",x"A9",x"02",x"91",x"8E",x"D0", -- 0x05B0
    x"4C",x"A5",x"83",x"F0",x"11",x"B5",x"00",x"91", -- 0x05B8
    x"80",x"A9",x"02",x"91",x"8E",x"C8",x"91",x"8E", -- 0x05C0
    x"B5",x"04",x"91",x"80",x"D0",x"37",x"A5",x"85", -- 0x05C8
    x"C9",x"11",x"D0",x"11",x"B5",x"08",x"91",x"80", -- 0x05D0
    x"A9",x"02",x"91",x"8E",x"C8",x"91",x"8E",x"B5", -- 0x05D8
    x"0C",x"91",x"80",x"D0",x"20",x"B5",x"08",x"91", -- 0x05E0
    x"80",x"A9",x"02",x"91",x"8E",x"C8",x"91",x"8E", -- 0x05E8
    x"B5",x"0C",x"91",x"80",x"A0",x"16",x"B5",x"00", -- 0x05F0
    x"91",x"80",x"A9",x"02",x"91",x"8E",x"C8",x"91", -- 0x05F8
    x"8E",x"B5",x"04",x"91",x"80",x"A6",x"8B",x"CA", -- 0x0600
    x"30",x"2E",x"4C",x"5D",x"A5",x"86",x"82",x"B4", -- 0x0608
    x"38",x"B5",x"20",x"18",x"79",x"84",x"BC",x"C9", -- 0x0610
    x"40",x"B0",x"1E",x"85",x"84",x"B5",x"28",x"79", -- 0x0618
    x"88",x"BC",x"C9",x"70",x"B0",x"13",x"85",x"85", -- 0x0620
    x"20",x"84",x"A6",x"A5",x"84",x"4A",x"29",x"07", -- 0x0628
    x"AA",x"A0",x"00",x"B1",x"80",x"3D",x"4E",x"BB", -- 0x0630
    x"60",x"C9",x"00",x"60",x"A9",x"FF",x"8D",x"0A", -- 0x0638
    x"18",x"BD",x"9C",x"BC",x"D0",x"20",x"B5",x"20", -- 0x0640
    x"C5",x"90",x"D0",x"05",x"FE",x"9C",x"BC",x"D0", -- 0x0648
    x"15",x"B0",x"07",x"A9",x"01",x"8D",x"0A",x"18", -- 0x0650
    x"D0",x"0B",x"A5",x"90",x"D5",x"20",x"B0",x"05", -- 0x0658
    x"A9",x"03",x"8D",x"0A",x"18",x"60",x"B5",x"28", -- 0x0660
    x"C5",x"91",x"D0",x"05",x"DE",x"9C",x"BC",x"F0", -- 0x0668
    x"D5",x"B0",x"07",x"A9",x"02",x"8D",x"0A",x"18", -- 0x0670
    x"D0",x"09",x"A5",x"91",x"D5",x"28",x"B0",x"03", -- 0x0678
    x"EE",x"0A",x"18",x"60",x"AD",x"00",x"18",x"85", -- 0x0680
    x"80",x"AD",x"01",x"18",x"85",x"81",x"A5",x"85", -- 0x0688
    x"29",x"FE",x"0A",x"65",x"80",x"85",x"80",x"90", -- 0x0690
    x"02",x"E6",x"81",x"A5",x"84",x"4A",x"4A",x"4A", -- 0x0698
    x"4A",x"18",x"65",x"80",x"85",x"80",x"90",x"02", -- 0x06A0
    x"E6",x"81",x"60",x"AC",x"26",x"18",x"B9",x"C0", -- 0x06A8
    x"00",x"D5",x"20",x"F0",x"05",x"88",x"10",x"F6", -- 0x06B0
    x"30",x"09",x"B9",x"D0",x"00",x"D5",x"28",x"D0", -- 0x06B8
    x"F4",x"F0",x"37",x"AC",x"09",x"18",x"30",x"17", -- 0x06C0
    x"B9",x"50",x"00",x"D5",x"20",x"F0",x"05",x"88", -- 0x06C8
    x"10",x"F4",x"30",x"0B",x"B9",x"5F",x"00",x"D5", -- 0x06D0
    x"28",x"D0",x"F4",x"A9",x"0F",x"D0",x"1D",x"86", -- 0x06D8
    x"8B",x"A4",x"7F",x"B9",x"20",x"00",x"D5",x"20", -- 0x06E0
    x"F0",x"05",x"88",x"10",x"F6",x"30",x"0F",x"C4", -- 0x06E8
    x"8B",x"F0",x"F7",x"B9",x"28",x"00",x"D5",x"28", -- 0x06F0
    x"D0",x"F0",x"A9",x"07",x"95",x"48",x"60",x"80", -- 0x06F8
    x"A0",x"C0",x"E0",x"00",x"20",x"40",x"16",x"16", -- 0x0700
    x"16",x"16",x"17",x"17",x"17",x"3F",x"CF",x"F3", -- 0x0708
    x"FC",x"00",x"00",x"00",x"00",x"40",x"10",x"04", -- 0x0710
    x"01",x"C0",x"30",x"0C",x"03",x"A0",x"E0",x"A9", -- 0x0718
    x"AA",x"99",x"7F",x"16",x"88",x"D0",x"FA",x"A9", -- 0x0720
    x"19",x"85",x"8E",x"A9",x"A7",x"85",x"8F",x"AE", -- 0x0728
    x"21",x"18",x"BD",x"0D",x"18",x"85",x"86",x"BD", -- 0x0730
    x"17",x"18",x"85",x"87",x"20",x"72",x"A7",x"CA", -- 0x0738
    x"D0",x"06",x"AD",x"22",x"18",x"F0",x"01",x"CA", -- 0x0740
    x"10",x"E8",x"A9",x"15",x"85",x"8E",x"A9",x"A7", -- 0x0748
    x"85",x"8F",x"A6",x"7F",x"B5",x"20",x"85",x"86", -- 0x0750
    x"B5",x"28",x"85",x"87",x"20",x"72",x"A7",x"CA", -- 0x0758
    x"10",x"F2",x"A9",x"11",x"85",x"8E",x"A9",x"A7", -- 0x0760
    x"85",x"8F",x"A5",x"90",x"85",x"86",x"A5",x"91", -- 0x0768
    x"85",x"87",x"A5",x"87",x"4A",x"4A",x"4A",x"4A", -- 0x0770
    x"A8",x"A5",x"86",x"29",x"F0",x"4A",x"79",x"FF", -- 0x0778
    x"A6",x"85",x"80",x"B9",x"06",x"A7",x"69",x"00", -- 0x0780
    x"85",x"81",x"A5",x"86",x"4A",x"4A",x"29",x"03", -- 0x0788
    x"85",x"89",x"A5",x"87",x"4A",x"29",x"06",x"A8", -- 0x0790
    x"85",x"8A",x"B1",x"80",x"A4",x"89",x"39",x"0D", -- 0x0798
    x"A7",x"11",x"8E",x"A4",x"8A",x"91",x"80",x"C8", -- 0x07A0
    x"91",x"80",x"60",x"AD",x"00",x"18",x"85",x"80", -- 0x07A8
    x"AD",x"01",x"18",x"85",x"81",x"A2",x"00",x"86", -- 0x07B0
    x"86",x"A5",x"91",x"4A",x"38",x"E9",x"04",x"85", -- 0x07B8
    x"87",x"10",x"17",x"8A",x"38",x"E5",x"87",x"85", -- 0x07C0
    x"87",x"0A",x"0A",x"85",x"86",x"A5",x"80",x"38", -- 0x07C8
    x"E5",x"86",x"85",x"80",x"B0",x"02",x"C6",x"81", -- 0x07D0
    x"D0",x"10",x"0A",x"26",x"86",x"0A",x"26",x"86", -- 0x07D8
    x"65",x"80",x"85",x"80",x"A5",x"86",x"65",x"81", -- 0x07E0
    x"85",x"81",x"A5",x"90",x"4A",x"38",x"E9",x"04", -- 0x07E8
    x"10",x"0D",x"A5",x"80",x"38",x"E9",x"01",x"85", -- 0x07F0
    x"80",x"A9",x"00",x"B0",x"02",x"C6",x"81",x"4A", -- 0x07F8
    x"4A",x"4A",x"18",x"65",x"80",x"85",x"80",x"90", -- 0x0800
    x"02",x"E6",x"81",x"A5",x"91",x"4A",x"38",x"E9", -- 0x0808
    x"04",x"8D",x"07",x"18",x"A9",x"6E",x"85",x"82", -- 0x0810
    x"A9",x"1E",x"85",x"83",x"A9",x"84",x"85",x"84", -- 0x0818
    x"A9",x"1E",x"85",x"85",x"A9",x"6E",x"85",x"8E", -- 0x0820
    x"A9",x"96",x"85",x"8F",x"A9",x"84",x"85",x"EB", -- 0x0828
    x"A9",x"96",x"85",x"EC",x"A5",x"91",x"4A",x"B0", -- 0x0830
    x"22",x"A5",x"90",x"4A",x"90",x"00",x"90",x"03", -- 0x0838
    x"4C",x"C6",x"A8",x"A9",x"09",x"85",x"88",x"0A", -- 0x0840
    x"8D",x"08",x"18",x"20",x"45",x"A9",x"20",x"0D", -- 0x0848
    x"A9",x"EE",x"07",x"18",x"C6",x"88",x"D0",x"F3", -- 0x0850
    x"4C",x"BC",x"A9",x"A9",x"6E",x"85",x"84",x"A9", -- 0x0858
    x"1E",x"85",x"85",x"A9",x"6E",x"85",x"EB",x"A9", -- 0x0860
    x"96",x"85",x"EC",x"A9",x"12",x"8D",x"08",x"18", -- 0x0868
    x"20",x"45",x"A9",x"20",x"0D",x"A9",x"EE",x"07", -- 0x0870
    x"18",x"A9",x"84",x"85",x"82",x"A9",x"1E",x"85", -- 0x0878
    x"83",x"A9",x"9A",x"85",x"84",x"A9",x"1E",x"85", -- 0x0880
    x"85",x"A9",x"84",x"85",x"8E",x"A9",x"96",x"85", -- 0x0888
    x"8F",x"A9",x"9A",x"85",x"EB",x"A9",x"96",x"85", -- 0x0890
    x"EC",x"A9",x"08",x"85",x"88",x"20",x"45",x"A9", -- 0x0898
    x"20",x"0D",x"A9",x"EE",x"07",x"18",x"C6",x"88", -- 0x08A0
    x"D0",x"F3",x"A5",x"84",x"38",x"E9",x"16",x"85", -- 0x08A8
    x"84",x"B0",x"02",x"C6",x"85",x"A5",x"EB",x"38", -- 0x08B0
    x"E9",x"16",x"85",x"EB",x"B0",x"02",x"C6",x"EC", -- 0x08B8
    x"20",x"45",x"A9",x"4C",x"BC",x"A9",x"A9",x"09", -- 0x08C0
    x"85",x"88",x"A9",x"02",x"8D",x"08",x"18",x"20", -- 0x08C8
    x"45",x"A9",x"A2",x"10",x"E6",x"89",x"A5",x"86", -- 0x08D0
    x"18",x"69",x"08",x"85",x"86",x"A9",x"12",x"8D", -- 0x08D8
    x"08",x"18",x"20",x"51",x"A9",x"A9",x"11",x"8D", -- 0x08E0
    x"08",x"18",x"A2",x"01",x"C6",x"89",x"A5",x"86", -- 0x08E8
    x"38",x"E9",x"09",x"85",x"86",x"29",x"07",x"C9", -- 0x08F0
    x"07",x"D0",x"02",x"C6",x"89",x"20",x"51",x"A9", -- 0x08F8
    x"20",x"0D",x"A9",x"EE",x"07",x"18",x"C6",x"88", -- 0x0900
    x"D0",x"C0",x"4C",x"BC",x"A9",x"A5",x"80",x"18", -- 0x0908
    x"69",x"04",x"85",x"80",x"90",x"03",x"E6",x"81", -- 0x0910
    x"18",x"A5",x"82",x"69",x"2C",x"85",x"82",x"90", -- 0x0918
    x"03",x"E6",x"83",x"18",x"A5",x"84",x"69",x"2C", -- 0x0920
    x"85",x"84",x"90",x"03",x"E6",x"85",x"18",x"A5", -- 0x0928
    x"8E",x"69",x"2C",x"85",x"8E",x"90",x"03",x"E6", -- 0x0930
    x"8F",x"18",x"A5",x"EB",x"69",x"2C",x"85",x"EB", -- 0x0938
    x"90",x"02",x"E6",x"EC",x"60",x"A5",x"90",x"4A", -- 0x0940
    x"38",x"E9",x"04",x"85",x"86",x"A2",x"00",x"86", -- 0x0948
    x"89",x"AD",x"07",x"18",x"C9",x"38",x"B0",x"52", -- 0x0950
    x"8E",x"06",x"18",x"A5",x"86",x"C9",x"20",x"90", -- 0x0958
    x"04",x"A9",x"2A",x"D0",x"12",x"29",x"07",x"AA", -- 0x0960
    x"A4",x"89",x"B1",x"80",x"3D",x"4E",x"BB",x"D0", -- 0x0968
    x"04",x"A9",x"20",x"D0",x"02",x"A9",x"FF",x"AC", -- 0x0970
    x"06",x"18",x"91",x"82",x"91",x"84",x"C8",x"91", -- 0x0978
    x"82",x"91",x"84",x"C9",x"2A",x"F0",x"04",x"A9", -- 0x0980
    x"04",x"D0",x"02",x"A9",x"07",x"91",x"8E",x"91", -- 0x0988
    x"EB",x"88",x"91",x"8E",x"91",x"EB",x"C8",x"E6", -- 0x0990
    x"86",x"A5",x"86",x"29",x"07",x"D0",x"02",x"E6", -- 0x0998
    x"89",x"98",x"AA",x"E8",x"EC",x"08",x"18",x"D0", -- 0x09A0
    x"AF",x"60",x"A0",x"11",x"A9",x"2A",x"91",x"82", -- 0x09A8
    x"91",x"84",x"A9",x"07",x"91",x"8E",x"91",x"EB", -- 0x09B0
    x"88",x"10",x"F1",x"60",x"AE",x"26",x"18",x"B5", -- 0x09B8
    x"C0",x"85",x"8C",x"B5",x"D0",x"20",x"15",x"AB", -- 0x09C0
    x"D0",x"7C",x"A5",x"82",x"F0",x"12",x"A9",x"59", -- 0x09C8
    x"91",x"80",x"A9",x"00",x"91",x"8E",x"A0",x"16", -- 0x09D0
    x"91",x"8E",x"A9",x"5B",x"91",x"80",x"D0",x"66", -- 0x09D8
    x"A5",x"84",x"C9",x"11",x"D0",x"12",x"A9",x"58", -- 0x09E0
    x"91",x"80",x"A9",x"00",x"91",x"8E",x"A0",x"16", -- 0x09E8
    x"91",x"8E",x"A9",x"5A",x"91",x"80",x"D0",x"4E", -- 0x09F0
    x"A5",x"83",x"F0",x"11",x"A9",x"5A",x"91",x"80", -- 0x09F8
    x"A9",x"00",x"91",x"8E",x"C8",x"91",x"8E",x"A9", -- 0x0A00
    x"5B",x"91",x"80",x"D0",x"39",x"A5",x"85",x"C9", -- 0x0A08
    x"11",x"D0",x"11",x"A9",x"58",x"91",x"80",x"A9", -- 0x0A10
    x"00",x"91",x"8E",x"C8",x"91",x"8E",x"A9",x"59", -- 0x0A18
    x"91",x"80",x"D0",x"22",x"A0",x"00",x"A9",x"58", -- 0x0A20
    x"91",x"80",x"A9",x"00",x"91",x"8E",x"C8",x"91", -- 0x0A28
    x"8E",x"A9",x"59",x"91",x"80",x"A0",x"16",x"A9", -- 0x0A30
    x"5A",x"91",x"80",x"A9",x"00",x"91",x"8E",x"C8", -- 0x0A38
    x"91",x"8E",x"A9",x"5B",x"91",x"80",x"CA",x"30", -- 0x0A40
    x"03",x"4C",x"BF",x"A9",x"AE",x"21",x"18",x"BD", -- 0x0A48
    x"0D",x"18",x"85",x"8C",x"BD",x"17",x"18",x"20", -- 0x0A50
    x"15",x"AB",x"D0",x"76",x"A5",x"82",x"F0",x"10", -- 0x0A58
    x"A9",x"51",x"91",x"80",x"A9",x"07",x"91",x"8E", -- 0x0A60
    x"A0",x"16",x"A9",x"20",x"91",x"80",x"D0",x"62", -- 0x0A68
    x"A5",x"84",x"C9",x"11",x"D0",x"12",x"A9",x"50", -- 0x0A70
    x"91",x"80",x"A9",x"07",x"91",x"8E",x"A0",x"16", -- 0x0A78
    x"91",x"8E",x"A9",x"52",x"91",x"80",x"D0",x"4A", -- 0x0A80
    x"A5",x"83",x"F0",x"0F",x"A9",x"52",x"91",x"80", -- 0x0A88
    x"A9",x"07",x"91",x"8E",x"C8",x"A9",x"20",x"91", -- 0x0A90
    x"80",x"D0",x"37",x"A5",x"85",x"C9",x"11",x"D0", -- 0x0A98
    x"11",x"A9",x"50",x"91",x"80",x"A9",x"07",x"91", -- 0x0AA0
    x"8E",x"C8",x"91",x"8E",x"A9",x"51",x"91",x"80", -- 0x0AA8
    x"D0",x"20",x"A0",x"00",x"A9",x"50",x"91",x"80", -- 0x0AB0
    x"A9",x"07",x"91",x"8E",x"C8",x"91",x"8E",x"A9", -- 0x0AB8
    x"51",x"91",x"80",x"A0",x"16",x"A9",x"52",x"91", -- 0x0AC0
    x"80",x"A9",x"07",x"91",x"8E",x"C8",x"A9",x"20", -- 0x0AC8
    x"91",x"80",x"CA",x"D0",x"06",x"AD",x"22",x"18", -- 0x0AD0
    x"F0",x"01",x"CA",x"30",x"03",x"4C",x"4F",x"AA", -- 0x0AD8
    x"98",x"30",x"27",x"A0",x"17",x"AD",x"22",x"18", -- 0x0AE0
    x"D0",x"20",x"A5",x"83",x"F0",x"02",x"A0",x"01", -- 0x0AE8
    x"A5",x"82",x"F0",x"02",x"A0",x"16",x"A5",x"84", -- 0x0AF0
    x"C9",x"11",x"F0",x"0E",x"A5",x"85",x"C9",x"11", -- 0x0AF8
    x"F0",x"08",x"A9",x"53",x"91",x"80",x"A9",x"02", -- 0x0B00
    x"91",x"8E",x"AD",x"0B",x"18",x"C9",x"09",x"90", -- 0x0B08
    x"03",x"4C",x"5B",x"A5",x"60",x"A0",x"00",x"84", -- 0x0B10
    x"82",x"84",x"83",x"38",x"E5",x"91",x"18",x"69", -- 0x0B18
    x"08",x"85",x"85",x"C9",x"12",x"90",x"08",x"C9", -- 0x0B20
    x"FF",x"D0",x"33",x"85",x"83",x"84",x"85",x"A5", -- 0x0B28
    x"8C",x"38",x"E5",x"90",x"18",x"69",x"08",x"85", -- 0x0B30
    x"84",x"C9",x"12",x"90",x"0A",x"C9",x"FF",x"D0", -- 0x0B38
    x"1D",x"85",x"82",x"84",x"84",x"98",x"18",x"A4", -- 0x0B40
    x"85",x"79",x"18",x"BB",x"85",x"80",x"85",x"8E", -- 0x0B48
    x"B9",x"2A",x"BB",x"69",x"00",x"85",x"81",x"49", -- 0x0B50
    x"88",x"85",x"8F",x"A0",x"00",x"60",x"A0",x"FF", -- 0x0B58
    x"60",x"EA",x"EA",x"A0",x"00",x"60",x"A0",x"FF", -- 0x0B60
    x"60",x"A9",x"00",x"85",x"95",x"A5",x"93",x"4A", -- 0x0B68
    x"90",x"03",x"4C",x"E7",x"AB",x"AD",x"3F",x"18", -- 0x0B70
    x"D0",x"05",x"20",x"C3",x"B1",x"D0",x"03",x"20", -- 0x0B78
    x"2E",x"A4",x"A5",x"E3",x"30",x"32",x"C5",x"8D", -- 0x0B80
    x"F0",x"2E",x"A6",x"E3",x"20",x"5A",x"AC",x"C9", -- 0x0B88
    x"FF",x"F0",x"25",x"C9",x"2A",x"F0",x"21",x"A5", -- 0x0B90
    x"8D",x"85",x"86",x"A5",x"E3",x"85",x"8D",x"38", -- 0x0B98
    x"E5",x"86",x"29",x"03",x"C9",x"02",x"F0",x"04", -- 0x0BA0
    x"E6",x"95",x"D0",x"56",x"A5",x"8D",x"38",x"E9", -- 0x0BA8
    x"01",x"29",x"03",x"85",x"92",x"4C",x"06",x"AC", -- 0x0BB0
    x"A6",x"8D",x"20",x"5A",x"AC",x"C9",x"FF",x"F0", -- 0x0BB8
    x"04",x"C9",x"2A",x"D0",x"22",x"E6",x"95",x"E6", -- 0x0BC0
    x"8D",x"A5",x"8D",x"29",x"03",x"85",x"8D",x"AA", -- 0x0BC8
    x"20",x"5A",x"AC",x"C9",x"FF",x"F0",x"04",x"C9", -- 0x0BD0
    x"2A",x"D0",x"27",x"E6",x"8D",x"E6",x"8D",x"A5", -- 0x0BD8
    x"8D",x"29",x"03",x"85",x"8D",x"10",x"1B",x"A4", -- 0x0BE0
    x"8D",x"B8",x"D0",x"04",x"C6",x"91",x"50",x"10", -- 0x0BE8
    x"88",x"D0",x"04",x"E6",x"90",x"50",x"09",x"88", -- 0x0BF0
    x"D0",x"04",x"E6",x"91",x"50",x"02",x"C6",x"90", -- 0x0BF8
    x"E6",x"93",x"A5",x"8D",x"85",x"92",x"20",x"AB", -- 0x0C00
    x"A7",x"A9",x"26",x"85",x"80",x"A9",x"1F",x"85", -- 0x0C08
    x"81",x"A9",x"26",x"85",x"8E",x"A9",x"97",x"85", -- 0x0C10
    x"8F",x"A2",x"01",x"BC",x"45",x"BC",x"B1",x"80", -- 0x0C18
    x"C9",x"50",x"90",x"0F",x"C9",x"55",x"B0",x"0B", -- 0x0C20
    x"A5",x"93",x"4A",x"B0",x"06",x"20",x"D8",x"B5", -- 0x0C28
    x"4C",x"36",x"AC",x"CA",x"10",x"E5",x"20",x"AF", -- 0x0C30
    x"AC",x"A5",x"92",x"D0",x"05",x"20",x"69",x"AC", -- 0x0C38
    x"30",x"15",x"C9",x"01",x"D0",x"05",x"20",x"77", -- 0x0C40
    x"AC",x"30",x"0C",x"C9",x"02",x"D0",x"05",x"20", -- 0x0C48
    x"85",x"AC",x"30",x"03",x"20",x"93",x"AC",x"4C", -- 0x0C50
    x"BE",x"AC",x"A0",x"00",x"BD",x"5C",x"BC",x"85", -- 0x0C58
    x"80",x"BD",x"60",x"BC",x"85",x"81",x"B1",x"80", -- 0x0C60
    x"60",x"A2",x"03",x"BC",x"44",x"BC",x"BD",x"48", -- 0x0C68
    x"BC",x"91",x"80",x"CA",x"10",x"F5",x"60",x"A2", -- 0x0C70
    x"03",x"BC",x"44",x"BC",x"BD",x"4C",x"BC",x"91", -- 0x0C78
    x"80",x"CA",x"10",x"F5",x"60",x"A2",x"03",x"BC", -- 0x0C80
    x"44",x"BC",x"BD",x"50",x"BC",x"91",x"80",x"CA", -- 0x0C88
    x"10",x"F5",x"60",x"A2",x"03",x"BC",x"44",x"BC", -- 0x0C90
    x"BD",x"54",x"BC",x"91",x"80",x"CA",x"10",x"F5", -- 0x0C98
    x"60",x"A2",x"03",x"BC",x"44",x"BC",x"BD",x"58", -- 0x0CA0
    x"BC",x"91",x"80",x"CA",x"10",x"F5",x"60",x"A9", -- 0x0CA8
    x"06",x"8D",x"26",x"97",x"8D",x"27",x"97",x"8D", -- 0x0CB0
    x"3C",x"97",x"8D",x"3D",x"97",x"60",x"A5",x"93", -- 0x0CB8
    x"4A",x"90",x"03",x"4C",x"45",x"AD",x"A5",x"95", -- 0x0CC0
    x"D0",x"7B",x"A5",x"7E",x"C9",x"04",x"F0",x"75", -- 0x0CC8
    x"A5",x"E2",x"F0",x"71",x"A5",x"8D",x"18",x"69", -- 0x0CD0
    x"02",x"29",x"03",x"85",x"8B",x"AA",x"20",x"5A", -- 0x0CD8
    x"AC",x"C9",x"2A",x"F0",x"60",x"C9",x"FF",x"F0", -- 0x0CE0
    x"5C",x"A5",x"94",x"D0",x"08",x"A5",x"E4",x"F0", -- 0x0CE8
    x"54",x"A9",x"03",x"85",x"94",x"20",x"70",x"B6", -- 0x0CF0
    x"A0",x"0E",x"88",x"30",x"1C",x"B9",x"50",x"00", -- 0x0CF8
    x"48",x"B9",x"5F",x"00",x"48",x"B9",x"6E",x"00", -- 0x0D00
    x"48",x"C8",x"68",x"99",x"6E",x"00",x"68",x"99", -- 0x0D08
    x"5F",x"00",x"68",x"99",x"50",x"00",x"88",x"10", -- 0x0D10
    x"E1",x"A4",x"8B",x"A5",x"90",x"18",x"79",x"84", -- 0x0D18
    x"BC",x"85",x"50",x"A5",x"91",x"18",x"79",x"88", -- 0x0D20
    x"BC",x"85",x"5F",x"A9",x"32",x"85",x"6E",x"AD", -- 0x0D28
    x"09",x"18",x"C9",x"0E",x"F0",x"05",x"EE",x"09", -- 0x0D30
    x"18",x"69",x"01",x"C6",x"94",x"EE",x"3B",x"18", -- 0x0D38
    x"A9",x"F2",x"8D",x"0B",x"90",x"AE",x"09",x"18", -- 0x0D40
    x"30",x"0C",x"B5",x"6E",x"D0",x"03",x"CE",x"09", -- 0x0D48
    x"18",x"D6",x"6E",x"CA",x"10",x"FB",x"AE",x"09", -- 0x0D50
    x"18",x"10",x"03",x"60",x"EA",x"EA",x"B5",x"50", -- 0x0D58
    x"85",x"8C",x"B5",x"5F",x"20",x"15",x"AB",x"D0", -- 0x0D60
    x"7C",x"A5",x"82",x"F0",x"12",x"A9",x"55",x"91", -- 0x0D68
    x"80",x"A9",x"01",x"91",x"8E",x"A0",x"16",x"91", -- 0x0D70
    x"8E",x"A9",x"57",x"91",x"80",x"D0",x"66",x"A5", -- 0x0D78
    x"84",x"C9",x"11",x"D0",x"12",x"A9",x"54",x"91", -- 0x0D80
    x"80",x"A9",x"01",x"91",x"8E",x"A0",x"16",x"91", -- 0x0D88
    x"8E",x"A9",x"56",x"91",x"80",x"D0",x"4E",x"A5", -- 0x0D90
    x"83",x"F0",x"11",x"A9",x"56",x"91",x"80",x"A9", -- 0x0D98
    x"01",x"91",x"8E",x"C8",x"91",x"8E",x"A9",x"57", -- 0x0DA0
    x"91",x"80",x"D0",x"39",x"A5",x"85",x"C9",x"11", -- 0x0DA8
    x"D0",x"11",x"A9",x"54",x"91",x"80",x"A9",x"01", -- 0x0DB0
    x"91",x"8E",x"C8",x"91",x"8E",x"A9",x"55",x"91", -- 0x0DB8
    x"80",x"D0",x"22",x"A0",x"00",x"A9",x"54",x"91", -- 0x0DC0
    x"80",x"A9",x"01",x"91",x"8E",x"C8",x"91",x"8E", -- 0x0DC8
    x"A9",x"55",x"91",x"80",x"A0",x"16",x"A9",x"56", -- 0x0DD0
    x"91",x"80",x"A9",x"01",x"91",x"8E",x"C8",x"91", -- 0x0DD8
    x"8E",x"A9",x"57",x"91",x"80",x"CA",x"30",x"03", -- 0x0DE0
    x"4C",x"5E",x"AD",x"60",x"AD",x"24",x"18",x"30", -- 0x0DE8
    x"27",x"CE",x"24",x"18",x"D0",x"22",x"A9",x"14", -- 0x0DF0
    x"8D",x"24",x"18",x"EE",x"25",x"18",x"AD",x"25", -- 0x0DF8
    x"18",x"4A",x"B0",x"0A",x"A9",x"A0",x"8D",x"C4", -- 0x0E00
    x"1E",x"8D",x"C5",x"1E",x"D0",x"0A",x"A9",x"98", -- 0x0E08
    x"8D",x"C4",x"1E",x"A9",x"B2",x"8D",x"C5",x"1E", -- 0x0E10
    x"CE",x"30",x"18",x"D0",x"2C",x"A9",x"05",x"8D", -- 0x0E18
    x"30",x"18",x"AC",x"32",x"18",x"AD",x"31",x"18", -- 0x0E20
    x"C9",x"02",x"BE",x"F7",x"BC",x"B0",x"03",x"BE", -- 0x0E28
    x"07",x"BD",x"CE",x"32",x"18",x"10",x"0F",x"A9", -- 0x0E30
    x"0F",x"8D",x"32",x"18",x"CE",x"31",x"18",x"D0", -- 0x0E38
    x"05",x"A9",x"04",x"8D",x"31",x"18",x"8E",x"0B", -- 0x0E40
    x"90",x"CE",x"33",x"18",x"D0",x"13",x"A9",x"03", -- 0x0E48
    x"8D",x"33",x"18",x"AC",x"2F",x"18",x"30",x"09", -- 0x0E50
    x"B9",x"F3",x"BC",x"8D",x"0C",x"90",x"CE",x"2F", -- 0x0E58
    x"18",x"AC",x"34",x"18",x"30",x"09",x"B9",x"17", -- 0x0E60
    x"BD",x"8D",x"0C",x"90",x"CE",x"34",x"18",x"AD", -- 0x0E68
    x"3B",x"18",x"F0",x"0D",x"A5",x"9E",x"38",x"E9", -- 0x0E70
    x"03",x"D0",x"06",x"8D",x"0B",x"90",x"8D",x"3B", -- 0x0E78
    x"18",x"AD",x"2B",x"18",x"30",x"27",x"CE",x"2C", -- 0x0E80
    x"18",x"08",x"AD",x"2C",x"18",x"38",x"E9",x"05", -- 0x0E88
    x"D0",x"09",x"8D",x"0B",x"90",x"8D",x"0C",x"90", -- 0x0E90
    x"CE",x"2B",x"18",x"28",x"D0",x"0F",x"A9",x"18", -- 0x0E98
    x"8D",x"2C",x"18",x"A9",x"E4",x"8D",x"0B",x"90", -- 0x0EA0
    x"A9",x"C8",x"8D",x"0C",x"90",x"CE",x"2D",x"18", -- 0x0EA8
    x"D0",x"1B",x"A9",x"28",x"8D",x"2D",x"18",x"A5", -- 0x0EB0
    x"E2",x"D0",x"12",x"AD",x"0B",x"18",x"10",x"05", -- 0x0EB8
    x"A9",x"01",x"8D",x"0B",x"18",x"A5",x"7E",x"C9", -- 0x0EC0
    x"12",x"F0",x"02",x"E6",x"7E",x"AD",x"21",x"18", -- 0x0EC8
    x"D0",x"06",x"AD",x"22",x"18",x"F0",x"01",x"60", -- 0x0ED0
    x"4C",x"1D",x"A7",x"A9",x"14",x"85",x"86",x"A5", -- 0x0ED8
    x"7D",x"F0",x"FC",x"C6",x"7D",x"20",x"49",x"AE", -- 0x0EE0
    x"C6",x"86",x"D0",x"F3",x"A0",x"00",x"8C",x"0A", -- 0x0EE8
    x"90",x"8C",x"0B",x"90",x"8C",x"0C",x"90",x"A2", -- 0x0EF0
    x"0C",x"A5",x"7D",x"F0",x"FC",x"C6",x"7D",x"CA", -- 0x0EF8
    x"D0",x"F7",x"B9",x"EC",x"BC",x"8D",x"0C",x"90", -- 0x0F00
    x"C8",x"C0",x"07",x"D0",x"EA",x"A2",x"24",x"A5", -- 0x0F08
    x"7D",x"F0",x"FC",x"C6",x"7D",x"CA",x"D0",x"F7", -- 0x0F10
    x"8E",x"0C",x"90",x"A2",x"0C",x"A5",x"7D",x"F0", -- 0x0F18
    x"FC",x"C6",x"7D",x"CA",x"D0",x"F7",x"4C",x"AF", -- 0x0F20
    x"B6",x"20",x"29",x"A2",x"A9",x"2A",x"85",x"28", -- 0x0F28
    x"A9",x"13",x"8D",x"38",x"18",x"8D",x"36",x"18", -- 0x0F30
    x"8D",x"37",x"18",x"A9",x"0F",x"8D",x"39",x"18", -- 0x0F38
    x"A5",x"7D",x"F0",x"FC",x"C6",x"7D",x"CE",x"36", -- 0x0F40
    x"18",x"D0",x"3B",x"A9",x"03",x"8D",x"36",x"18", -- 0x0F48
    x"AD",x"38",x"18",x"30",x"31",x"20",x"5B",x"A5", -- 0x0F50
    x"C6",x"20",x"AC",x"38",x"18",x"C0",x"12",x"B0", -- 0x0F58
    x"0B",x"B9",x"7C",x"BB",x"99",x"F2",x"1E",x"A9", -- 0x0F60
    x"20",x"99",x"DC",x"1E",x"CE",x"38",x"18",x"D0", -- 0x0F68
    x"15",x"A0",x"02",x"B9",x"90",x"BB",x"99",x"25", -- 0x0F70
    x"1F",x"88",x"10",x"F7",x"AD",x"35",x"18",x"29", -- 0x0F78
    x"0F",x"09",x"30",x"8D",x"28",x"1F",x"CE",x"37", -- 0x0F80
    x"18",x"D0",x"B5",x"A9",x"0A",x"8D",x"37",x"18", -- 0x0F88
    x"AC",x"39",x"18",x"B9",x"38",x"BD",x"8D",x"0C", -- 0x0F90
    x"90",x"CE",x"39",x"18",x"10",x"A2",x"EE",x"35", -- 0x0F98
    x"18",x"A9",x"CE",x"8D",x"0F",x"90",x"60",x"20", -- 0x0FA0
    x"E6",x"AF",x"20",x"CD",x"B8",x"A9",x"00",x"8D", -- 0x0FA8
    x"0A",x"90",x"8D",x"0B",x"90",x"8D",x"0C",x"90", -- 0x0FB0
    x"A9",x"7F",x"8D",x"0E",x"90",x"A0",x"2E",x"A5", -- 0x0FB8
    x"7D",x"F0",x"FC",x"C6",x"7D",x"CE",x"2E",x"18", -- 0x0FC0
    x"D0",x"F5",x"A9",x"06",x"8D",x"2E",x"18",x"B9", -- 0x0FC8
    x"48",x"BD",x"8D",x"0C",x"90",x"C0",x"12",x"D0", -- 0x0FD0
    x"07",x"98",x"48",x"20",x"00",x"B0",x"68",x"A8", -- 0x0FD8
    x"88",x"10",x"DC",x"4C",x"A4",x"B7",x"A2",x"03", -- 0x0FE0
    x"86",x"9F",x"A2",x"01",x"86",x"E0",x"8E",x"35", -- 0x0FE8
    x"18",x"CA",x"86",x"E5",x"86",x"E7",x"86",x"E9", -- 0x0FF0
    x"86",x"9C",x"8E",x"3C",x"18",x"86",x"E1",x"60", -- 0x0FF8
    x"A9",x"00",x"85",x"80",x"A9",x"1E",x"85",x"81", -- 0x1000
    x"A9",x"00",x"85",x"8E",x"A9",x"96",x"85",x"8F", -- 0x1008
    x"A2",x"04",x"A0",x"00",x"A9",x"A0",x"91",x"80", -- 0x1010
    x"A9",x"06",x"91",x"8E",x"88",x"D0",x"F5",x"E6", -- 0x1018
    x"81",x"E6",x"8F",x"CA",x"D0",x"EC",x"A0",x"88", -- 0x1020
    x"8C",x"0D",x"1E",x"C8",x"8C",x"0E",x"1E",x"A0", -- 0x1028
    x"04",x"B9",x"56",x"BB",x"99",x"01",x"1E",x"88", -- 0x1030
    x"10",x"F7",x"A0",x"0D",x"B9",x"5B",x"BB",x"99", -- 0x1038
    x"2D",x"1E",x"88",x"10",x"F7",x"A9",x"00",x"20", -- 0x1040
    x"BA",x"B1",x"A2",x"07",x"BC",x"93",x"BB",x"BD", -- 0x1048
    x"69",x"BB",x"99",x"80",x"1E",x"CA",x"10",x"F4", -- 0x1050
    x"A9",x"B0",x"8D",x"AE",x"1E",x"8D",x"AF",x"1E", -- 0x1058
    x"A0",x"02",x"B9",x"71",x"BB",x"99",x"EE",x"1E", -- 0x1060
    x"88",x"10",x"F7",x"A5",x"E0",x"29",x"0F",x"09", -- 0x1068
    x"B0",x"8D",x"07",x"1F",x"A5",x"E0",x"4A",x"4A", -- 0x1070
    x"4A",x"4A",x"F0",x"05",x"09",x"B0",x"8D",x"06", -- 0x1078
    x"1F",x"A9",x"30",x"85",x"80",x"A9",x"1F",x"85", -- 0x1080
    x"81",x"A9",x"30",x"85",x"8E",x"A9",x"97",x"85", -- 0x1088
    x"8F",x"A2",x"D0",x"A9",x"06",x"85",x"86",x"A0", -- 0x1090
    x"00",x"A9",x"08",x"91",x"8E",x"8A",x"91",x"80", -- 0x1098
    x"E8",x"C8",x"C0",x"04",x"D0",x"F3",x"A5",x"80", -- 0x10A0
    x"69",x"15",x"85",x"80",x"85",x"8E",x"90",x"04", -- 0x10A8
    x"E6",x"81",x"E6",x"8F",x"C6",x"86",x"10",x"DF", -- 0x10B0
    x"A0",x"07",x"B9",x"8C",x"BC",x"99",x"20",x"00", -- 0x10B8
    x"B9",x"94",x"BC",x"99",x"28",x"00",x"A9",x"00", -- 0x10C0
    x"99",x"38",x"00",x"99",x"40",x"00",x"99",x"30", -- 0x10C8
    x"00",x"99",x"48",x"00",x"A9",x"20",x"99",x"4E", -- 0x10D0
    x"18",x"A9",x"EC",x"99",x"B0",x"00",x"A9",x"20", -- 0x10D8
    x"99",x"B8",x"00",x"88",x"10",x"D4",x"A9",x"1E", -- 0x10E0
    x"85",x"90",x"A9",x"64",x"85",x"91",x"20",x"AB", -- 0x10E8
    x"A7",x"A9",x"26",x"85",x"80",x"A9",x"1F",x"85", -- 0x10F0
    x"81",x"20",x"69",x"AC",x"20",x"AF",x"AC",x"20", -- 0x10F8
    x"5B",x"A5",x"A9",x"EC",x"85",x"96",x"A9",x"20", -- 0x1100
    x"85",x"97",x"A9",x"20",x"85",x"98",x"A2",x"01", -- 0x1108
    x"8E",x"30",x"18",x"8E",x"33",x"18",x"86",x"9E", -- 0x1110
    x"8E",x"2A",x"18",x"A2",x"04",x"8E",x"31",x"18", -- 0x1118
    x"A2",x"0F",x"8E",x"32",x"18",x"A2",x"50",x"86", -- 0x1120
    x"E2",x"CA",x"8E",x"0B",x"18",x"A4",x"E1",x"B9", -- 0x1128
    x"1E",x"BE",x"10",x"03",x"8D",x"0B",x"18",x"A2", -- 0x1130
    x"09",x"BD",x"0E",x"BB",x"9D",x"44",x"18",x"CA", -- 0x1138
    x"10",x"F7",x"86",x"9B",x"8E",x"24",x"18",x"8E", -- 0x1140
    x"2F",x"18",x"8E",x"34",x"18",x"8E",x"09",x"18", -- 0x1148
    x"8E",x"2B",x"18",x"E8",x"86",x"94",x"86",x"93", -- 0x1150
    x"86",x"8D",x"86",x"92",x"86",x"9D",x"8E",x"28", -- 0x1158
    x"18",x"8E",x"23",x"18",x"86",x"86",x"20",x"33", -- 0x1160
    x"B5",x"20",x"A1",x"B5",x"20",x"F4",x"B3",x"20", -- 0x1168
    x"1D",x"A7",x"4C",x"45",x"B6",x"A9",x"A0",x"85", -- 0x1170
    x"8B",x"A9",x"00",x"8D",x"27",x"18",x"A9",x"6E", -- 0x1178
    x"85",x"80",x"A9",x"1E",x"85",x"81",x"A2",x"11", -- 0x1180
    x"86",x"86",x"A9",x"6E",x"85",x"8E",x"A9",x"96", -- 0x1188
    x"85",x"8F",x"A4",x"86",x"A5",x"8B",x"91",x"80", -- 0x1190
    x"AD",x"27",x"18",x"91",x"8E",x"88",x"10",x"F4", -- 0x1198
    x"A5",x"80",x"18",x"69",x"16",x"85",x"80",x"90", -- 0x11A0
    x"02",x"E6",x"81",x"A5",x"8E",x"18",x"69",x"16", -- 0x11A8
    x"85",x"8E",x"90",x"02",x"E6",x"8F",x"CA",x"10", -- 0x11B0
    x"D9",x"60",x"A0",x"09",x"99",x"31",x"96",x"88", -- 0x11B8
    x"10",x"FA",x"60",x"A2",x"00",x"86",x"E4",x"A2", -- 0x11C0
    x"03",x"BD",x"3C",x"BB",x"8D",x"20",x"91",x"AD", -- 0x11C8
    x"21",x"91",x"CD",x"21",x"91",x"D0",x"F8",x"3D", -- 0x11D0
    x"40",x"BB",x"F0",x"03",x"CA",x"10",x"EA",x"86", -- 0x11D8
    x"E3",x"A9",x"DF",x"8D",x"20",x"91",x"AD",x"21", -- 0x11E0
    x"91",x"CD",x"21",x"91",x"D0",x"F8",x"29",x"02", -- 0x11E8
    x"D0",x"02",x"E6",x"E4",x"78",x"A2",x"7F",x"8E", -- 0x11F0
    x"22",x"91",x"AD",x"20",x"91",x"CD",x"20",x"91", -- 0x11F8
    x"D0",x"F8",x"8E",x"20",x"91",x"A2",x"FF",x"8E", -- 0x1200
    x"22",x"91",x"58",x"29",x"80",x"D0",x"04",x"A9", -- 0x1208
    x"01",x"85",x"E3",x"AD",x"1F",x"91",x"CD",x"1F", -- 0x1210
    x"91",x"D0",x"F8",x"A8",x"A2",x"02",x"98",x"3D", -- 0x1218
    x"44",x"BB",x"D0",x"05",x"BD",x"47",x"BB",x"85", -- 0x1220
    x"E3",x"CA",x"10",x"F2",x"98",x"29",x"20",x"D0", -- 0x1228
    x"04",x"A9",x"01",x"85",x"E4",x"60",x"78",x"20", -- 0x1230
    x"8E",x"BA",x"F0",x"77",x"A2",x"02",x"BD",x"BE", -- 0x1238
    x"B2",x"8D",x"20",x"91",x"AD",x"21",x"91",x"CD", -- 0x1240
    x"21",x"91",x"D0",x"F8",x"3D",x"C1",x"B2",x"D0", -- 0x1248
    x"06",x"CA",x"10",x"EA",x"8E",x"43",x"18",x"CE", -- 0x1250
    x"40",x"18",x"D0",x"57",x"A9",x"04",x"8D",x"40", -- 0x1258
    x"18",x"A2",x"03",x"BD",x"4A",x"BB",x"8D",x"20", -- 0x1260
    x"91",x"AD",x"21",x"91",x"10",x"05",x"CA",x"10", -- 0x1268
    x"F2",x"30",x"1F",x"18",x"8A",x"F0",x"27",x"CA", -- 0x1270
    x"F0",x"2F",x"CA",x"F0",x"0B",x"8A",x"6D",x"01", -- 0x1278
    x"90",x"29",x"3F",x"8D",x"01",x"90",x"90",x"0A", -- 0x1280
    x"AD",x"00",x"90",x"69",x"01",x"29",x"8F",x"8D", -- 0x1288
    x"00",x"90",x"AD",x"1F",x"91",x"CD",x"1F",x"91", -- 0x1290
    x"D0",x"F8",x"29",x"20",x"D0",x"15",x"A2",x"FA", -- 0x1298
    x"9A",x"CE",x"3F",x"18",x"D8",x"58",x"4C",x"1E", -- 0x12A0
    x"B4",x"AD",x"00",x"90",x"49",x"80",x"8D",x"00", -- 0x12A8
    x"90",x"90",x"DF",x"68",x"A8",x"68",x"AA",x"68", -- 0x12B0
    x"40",x"EA",x"EA",x"EA",x"EA",x"EA",x"F7",x"EF", -- 0x12B8
    x"DF",x"02",x"40",x"01",x"A2",x"50",x"A5",x"7D", -- 0x12C0
    x"F0",x"FC",x"C6",x"7D",x"CA",x"D0",x"F7",x"60", -- 0x12C8
    x"A2",x"0B",x"0E",x"3D",x"18",x"2E",x"3E",x"18", -- 0x12D0
    x"2A",x"2A",x"4D",x"3D",x"18",x"2A",x"4D",x"3D", -- 0x12D8
    x"18",x"4A",x"4A",x"49",x"FF",x"29",x"01",x"0D", -- 0x12E0
    x"3D",x"18",x"8D",x"3D",x"18",x"CA",x"D0",x"E2", -- 0x12E8
    x"38",x"E5",x"8B",x"C5",x"8B",x"B0",x"F9",x"0A", -- 0x12F0
    x"60",x"AD",x"02",x"18",x"85",x"80",x"AD",x"03", -- 0x12F8
    x"18",x"85",x"81",x"AD",x"04",x"18",x"85",x"82", -- 0x1300
    x"AD",x"05",x"18",x"85",x"83",x"A0",x"0F",x"B1", -- 0x1308
    x"80",x"99",x"C0",x"00",x"B1",x"82",x"99",x"D0", -- 0x1310
    x"00",x"88",x"10",x"F3",x"A4",x"E1",x"B9",x"1E", -- 0x1318
    x"BE",x"30",x"2B",x"A9",x"10",x"85",x"8B",x"A2", -- 0x1320
    x"07",x"8A",x"48",x"20",x"D0",x"B2",x"4A",x"A8", -- 0x1328
    x"C8",x"C0",x"10",x"F0",x"12",x"B9",x"C0",x"00", -- 0x1330
    x"48",x"B9",x"D0",x"00",x"88",x"99",x"D0",x"00", -- 0x1338
    x"68",x"99",x"C0",x"00",x"C8",x"10",x"E9",x"C6", -- 0x1340
    x"8B",x"68",x"AA",x"CA",x"10",x"DB",x"A2",x"09", -- 0x1348
    x"8A",x"48",x"A9",x"20",x"85",x"8B",x"20",x"D0", -- 0x1350
    x"B2",x"85",x"84",x"A9",x"38",x"85",x"8B",x"20", -- 0x1358
    x"D0",x"B2",x"85",x"85",x"20",x"84",x"A6",x"A0", -- 0x1360
    x"00",x"A5",x"84",x"4A",x"29",x"07",x"AA",x"B1", -- 0x1368
    x"80",x"3D",x"4E",x"BB",x"D0",x"DC",x"68",x"AA", -- 0x1370
    x"A8",x"A5",x"84",x"4A",x"4A",x"4A",x"85",x"8A", -- 0x1378
    x"C8",x"C0",x"0A",x"F0",x"1F",x"B9",x"0D",x"18", -- 0x1380
    x"4A",x"4A",x"4A",x"C5",x"8A",x"D0",x"F1",x"B9", -- 0x1388
    x"17",x"18",x"4A",x"4A",x"4A",x"85",x"8A",x"A5", -- 0x1390
    x"85",x"4A",x"4A",x"4A",x"C5",x"8A",x"D0",x"D9", -- 0x1398
    x"8A",x"48",x"10",x"AE",x"A0",x"0F",x"A5",x"84", -- 0x13A0
    x"D9",x"C0",x"00",x"F0",x"05",x"88",x"10",x"F6", -- 0x13A8
    x"30",x"09",x"A5",x"85",x"D9",x"D0",x"00",x"D0", -- 0x13B0
    x"F4",x"F0",x"E5",x"A0",x"07",x"A5",x"84",x"4A", -- 0x13B8
    x"4A",x"4A",x"85",x"8A",x"88",x"30",x"1D",x"B9", -- 0x13C0
    x"8C",x"BC",x"4A",x"4A",x"4A",x"C5",x"8A",x"D0", -- 0x13C8
    x"F3",x"B9",x"94",x"BC",x"4A",x"4A",x"4A",x"85", -- 0x13D0
    x"8A",x"A5",x"85",x"4A",x"4A",x"4A",x"C5",x"8A", -- 0x13D8
    x"D0",x"DB",x"F0",x"BC",x"A5",x"84",x"9D",x"0D", -- 0x13E0
    x"18",x"A5",x"85",x"9D",x"17",x"18",x"CA",x"30", -- 0x13E8
    x"2C",x"4C",x"50",x"B3",x"A9",x"3C",x"85",x"80", -- 0x13F0
    x"A9",x"1E",x"85",x"81",x"A6",x"9F",x"CA",x"F0", -- 0x13F8
    x"1C",x"A0",x"00",x"A9",x"C0",x"91",x"80",x"C8", -- 0x1400
    x"A9",x"C1",x"91",x"80",x"A0",x"16",x"A9",x"C2", -- 0x1408
    x"91",x"80",x"C8",x"A9",x"C3",x"91",x"80",x"E6", -- 0x1410
    x"80",x"E6",x"80",x"D0",x"E1",x"60",x"20",x"75", -- 0x1418
    x"B1",x"A9",x"CE",x"8D",x"0F",x"90",x"AD",x"0E", -- 0x1420
    x"90",x"09",x"0F",x"8D",x"0E",x"90",x"A2",x"04", -- 0x1428
    x"A0",x"02",x"8C",x"0A",x"90",x"8C",x"0B",x"90", -- 0x1430
    x"A5",x"7D",x"F0",x"FC",x"C6",x"7D",x"88",x"D0", -- 0x1438
    x"F7",x"A0",x"02",x"A9",x"00",x"8D",x"0C",x"90", -- 0x1440
    x"BD",x"FA",x"B4",x"8D",x"0C",x"90",x"CA",x"10", -- 0x1448
    x"E7",x"A2",x"03",x"86",x"87",x"BD",x"9B",x"BB", -- 0x1450
    x"9D",x"9D",x"1E",x"CA",x"10",x"F7",x"A2",x"0B", -- 0x1458
    x"BD",x"9F",x"BB",x"9D",x"C8",x"1E",x"CA",x"10", -- 0x1460
    x"F7",x"A2",x"0D",x"BD",x"C5",x"BB",x"9D",x"37", -- 0x1468
    x"1F",x"CA",x"10",x"F7",x"A2",x"0C",x"BD",x"AB", -- 0x1470
    x"BB",x"9D",x"F5",x"1E",x"BD",x"B8",x"BB",x"9D", -- 0x1478
    x"0A",x"1F",x"CA",x"10",x"F1",x"A2",x"04",x"BD", -- 0x1480
    x"A6",x"BB",x"CA",x"10",x"FA",x"A2",x"0A",x"BC", -- 0x1488
    x"E9",x"BB",x"BD",x"D3",x"BB",x"99",x"A4",x"1F", -- 0x1490
    x"BD",x"DE",x"BB",x"99",x"C3",x"1F",x"CA",x"10", -- 0x1498
    x"EE",x"A9",x"13",x"8D",x"8D",x"1F",x"A9",x"10", -- 0x14A0
    x"8D",x"82",x"1F",x"A9",x"03",x"8D",x"35",x"1F", -- 0x14A8
    x"EA",x"A9",x"0C",x"8D",x"97",x"1F",x"A9",x"3B", -- 0x14B0
    x"8D",x"99",x"1F",x"A9",x"2E",x"8D",x"AE",x"1F", -- 0x14B8
    x"A2",x"11",x"A9",x"AD",x"9D",x"60",x"1F",x"CA", -- 0x14C0
    x"10",x"FA",x"A5",x"7D",x"F0",x"FC",x"C6",x"7D", -- 0x14C8
    x"20",x"A0",x"BA",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x14D0
    x"EA",x"EA",x"D0",x"03",x"4C",x"A7",x"AF",x"C6", -- 0x14D8
    x"87",x"D0",x"E7",x"A9",x"0A",x"85",x"87",x"E6", -- 0x14E0
    x"86",x"A5",x"86",x"4A",x"A9",x"02",x"90",x"02", -- 0x14E8
    x"A9",x"04",x"8D",x"9B",x"96",x"8D",x"A2",x"96", -- 0x14F0
    x"D0",x"D0",x"00",x"F3",x"F5",x"F4",x"F6",x"A2", -- 0x14F8
    x"00",x"BD",x"00",x"80",x"9D",x"00",x"10",x"BD", -- 0x1500
    x"00",x"81",x"9D",x"00",x"11",x"BD",x"0E",x"B9", -- 0x1508
    x"9D",x"00",x"12",x"49",x"FF",x"9D",x"00",x"16", -- 0x1510
    x"BD",x"0E",x"BA",x"9D",x"00",x"13",x"49",x"FF", -- 0x1518
    x"9D",x"00",x"17",x"BD",x"00",x"84",x"9D",x"00", -- 0x1520
    x"14",x"BD",x"00",x"85",x"9D",x"00",x"15",x"CA", -- 0x1528
    x"D0",x"CF",x"60",x"F8",x"A2",x"00",x"AD",x"3F", -- 0x1530
    x"18",x"D0",x"11",x"A5",x"86",x"18",x"65",x"E9", -- 0x1538
    x"85",x"E9",x"8A",x"65",x"E7",x"85",x"E7",x"8A", -- 0x1540
    x"65",x"E5",x"85",x"E5",x"D8",x"A5",x"E7",x"C9", -- 0x1548
    x"20",x"D0",x"17",x"A5",x"9C",x"D0",x"13",x"E6", -- 0x1550
    x"9F",x"E6",x"9C",x"A5",x"80",x"48",x"A5",x"81", -- 0x1558
    x"48",x"20",x"F4",x"B3",x"68",x"85",x"81",x"68", -- 0x1560
    x"85",x"80",x"A9",x"05",x"85",x"82",x"A9",x"1E", -- 0x1568
    x"85",x"83",x"A0",x"00",x"B9",x"E5",x"00",x"20", -- 0x1570
    x"BC",x"B5",x"C0",x"06",x"D0",x"F6",x"A9",x"B0", -- 0x1578
    x"91",x"82",x"A5",x"EA",x"C5",x"E9",x"A5",x"E8", -- 0x1580
    x"E5",x"E7",x"A5",x"E6",x"E5",x"E5",x"B0",x"2B", -- 0x1588
    x"A5",x"E5",x"85",x"E6",x"A5",x"E7",x"85",x"E8", -- 0x1590
    x"A5",x"E9",x"85",x"EA",x"A9",x"01",x"8D",x"3C", -- 0x1598
    x"18",x"A9",x"0E",x"85",x"82",x"A9",x"1E",x"85", -- 0x15A0
    x"83",x"A2",x"00",x"A0",x"00",x"B9",x"E6",x"00", -- 0x15A8
    x"20",x"BC",x"B5",x"C0",x"06",x"D0",x"F6",x"A9", -- 0x15B0
    x"B0",x"91",x"82",x"60",x"48",x"4A",x"4A",x"4A", -- 0x15B8
    x"4A",x"20",x"C7",x"B5",x"68",x"29",x"0F",x"D0", -- 0x15C0
    x"08",x"E0",x"00",x"D0",x"04",x"C0",x"05",x"D0", -- 0x15C8
    x"05",x"E8",x"09",x"B0",x"91",x"82",x"C8",x"60", -- 0x15D0
    x"AC",x"21",x"18",x"A5",x"91",x"D9",x"17",x"18", -- 0x15D8
    x"F0",x"03",x"88",x"10",x"F6",x"A5",x"90",x"D9", -- 0x15E0
    x"0D",x"18",x"D0",x"F6",x"EE",x"28",x"18",x"A9", -- 0x15E8
    x"03",x"8D",x"2F",x"18",x"84",x"9B",x"98",x"D0", -- 0x15F0
    x"12",x"A9",x"20",x"8D",x"34",x"18",x"A9",x"01", -- 0x15F8
    x"8D",x"24",x"18",x"8D",x"22",x"18",x"8D",x"23", -- 0x1600
    x"18",x"D0",x"22",x"AA",x"C8",x"C0",x"0A",x"F0", -- 0x1608
    x"0A",x"B9",x"0D",x"18",x"88",x"99",x"0D",x"18", -- 0x1610
    x"C8",x"10",x"F1",x"E8",x"E0",x"0A",x"F0",x"0A", -- 0x1618
    x"BD",x"17",x"18",x"CA",x"9D",x"17",x"18",x"E8", -- 0x1620
    x"10",x"F1",x"CE",x"21",x"18",x"AD",x"28",x"18", -- 0x1628
    x"0A",x"0A",x"0A",x"0A",x"C9",x"A0",x"F0",x"26", -- 0x1630
    x"85",x"86",x"20",x"33",x"B5",x"AD",x"23",x"18", -- 0x1638
    x"F0",x"03",x"20",x"33",x"B5",x"AD",x"28",x"18", -- 0x1640
    x"F8",x"18",x"69",x"01",x"AA",x"D8",x"29",x"10", -- 0x1648
    x"F0",x"05",x"A9",x"B1",x"8D",x"AC",x"1E",x"8A", -- 0x1650
    x"09",x"B0",x"8D",x"AD",x"1E",x"60",x"A9",x"50", -- 0x1658
    x"85",x"86",x"20",x"6A",x"B6",x"AD",x"23",x"18", -- 0x1660
    x"F0",x"F3",x"20",x"33",x"B5",x"4C",x"33",x"B5", -- 0x1668
    x"AD",x"3F",x"18",x"D0",x"E8",x"C6",x"E2",x"10", -- 0x1670
    x"02",x"E6",x"E2",x"A5",x"E2",x"C9",x"0C",x"D0", -- 0x1678
    x"19",x"A9",x"05",x"8D",x"2B",x"18",x"8D",x"2C", -- 0x1680
    x"18",x"AD",x"21",x"18",x"D0",x"05",x"AD",x"22", -- 0x1688
    x"18",x"D0",x"05",x"A9",x"02",x"20",x"BA",x"B1", -- 0x1690
    x"A5",x"E2",x"4A",x"4A",x"4A",x"A8",x"A5",x"E2", -- 0x1698
    x"29",x"07",x"D0",x"04",x"A9",x"A0",x"D0",x"03", -- 0x16A0
    x"18",x"69",x"77",x"99",x"31",x"1E",x"60",x"A2", -- 0x16A8
    x"00",x"86",x"7D",x"E8",x"85",x"86",x"A5",x"E2", -- 0x16B0
    x"D0",x"03",x"4C",x"C4",x"B2",x"A9",x"F0",x"8D", -- 0x16B8
    x"0C",x"90",x"20",x"70",x"B6",x"A9",x"06",x"85", -- 0x16C0
    x"87",x"A5",x"7D",x"F0",x"FC",x"C6",x"7D",x"20", -- 0x16C8
    x"33",x"B5",x"A5",x"87",x"38",x"E9",x"04",x"D0", -- 0x16D0
    x"03",x"8D",x"0C",x"90",x"C6",x"87",x"D0",x"E9", -- 0x16D8
    x"F0",x"D4",x"05",x"19",x"96",x"2E",x"00",x"FC", -- 0x16E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16E8
    x"70",x"5E",x"D8",x"78",x"A2",x"FF",x"9A",x"20", -- 0x16F0
    x"8A",x"FF",x"A2",x"0F",x"BD",x"E2",x"B6",x"9D", -- 0x16F8
    x"00",x"90",x"CA",x"10",x"F7",x"20",x"FF",x"B4", -- 0x1700
    x"A9",x"00",x"8D",x"1E",x"91",x"A9",x"C0",x"8D", -- 0x1708
    x"2E",x"91",x"A9",x"40",x"8D",x"1B",x"91",x"8D", -- 0x1710
    x"2B",x"91",x"A9",x"FF",x"8D",x"22",x"91",x"A9", -- 0x1718
    x"80",x"8D",x"13",x"91",x"A9",x"82",x"8D",x"1E", -- 0x1720
    x"91",x"A9",x"89",x"8D",x"24",x"91",x"A9",x"42", -- 0x1728
    x"8D",x"25",x"91",x"A9",x"36",x"8D",x"14",x"03", -- 0x1730
    x"A9",x"B2",x"8D",x"15",x"03",x"A0",x"1F",x"B9", -- 0x1738
    x"64",x"BC",x"99",x"00",x"00",x"88",x"10",x"F7", -- 0x1740
    x"C8",x"84",x"E6",x"84",x"EA",x"8C",x"3B",x"18", -- 0x1748
    x"8C",x"43",x"18",x"8C",x"3E",x"18",x"C8",x"8C", -- 0x1750
    x"2E",x"18",x"8C",x"3A",x"18",x"8C",x"3F",x"18", -- 0x1758
    x"8C",x"40",x"18",x"A9",x"4B",x"8D",x"3D",x"18", -- 0x1760
    x"A9",x"20",x"85",x"E8",x"EA",x"20",x"E6",x"AF", -- 0x1768
    x"20",x"CD",x"B8",x"A9",x"46",x"8D",x"29",x"18", -- 0x1770
    x"A2",x"06",x"A4",x"E1",x"B9",x"1E",x"BE",x"10", -- 0x1778
    x"10",x"A5",x"7F",x"48",x"20",x"29",x"AF",x"68", -- 0x1780
    x"85",x"7F",x"A9",x"23",x"8D",x"29",x"18",x"A2", -- 0x1788
    x"04",x"86",x"7E",x"AD",x"3A",x"18",x"F0",x"09", -- 0x1790
    x"20",x"00",x"B0",x"CE",x"3A",x"18",x"4C",x"C3", -- 0x1798
    x"A0",x"20",x"00",x"B0",x"20",x"C4",x"B2",x"20", -- 0x17A0
    x"1D",x"A7",x"A5",x"7D",x"F0",x"FC",x"C6",x"9E", -- 0x17A8
    x"D0",x"0E",x"A5",x"7E",x"85",x"9E",x"20",x"69", -- 0x17B0
    x"AB",x"20",x"A1",x"B8",x"A5",x"9D",x"D0",x"5B", -- 0x17B8
    x"AD",x"0B",x"18",x"30",x"10",x"CE",x"0B",x"18", -- 0x17C0
    x"D0",x"0B",x"A4",x"E1",x"B9",x"00",x"BE",x"8D", -- 0x17C8
    x"0B",x"18",x"20",x"7D",x"A4",x"CE",x"2A",x"18", -- 0x17D0
    x"D0",x"09",x"AD",x"29",x"18",x"8D",x"2A",x"18", -- 0x17D8
    x"20",x"70",x"B6",x"20",x"EC",x"AD",x"20",x"A1", -- 0x17E0
    x"B8",x"A5",x"9D",x"D0",x"2E",x"AD",x"21",x"18", -- 0x17E8
    x"D0",x"22",x"AD",x"22",x"18",x"F0",x"1D",x"20", -- 0x17F0
    x"5B",x"A5",x"20",x"DB",x"AE",x"E6",x"E1",x"A5", -- 0x17F8
    x"E1",x"38",x"E9",x"0F",x"D0",x"02",x"85",x"E1", -- 0x1800
    x"F8",x"A5",x"E0",x"18",x"69",x"01",x"85",x"E0", -- 0x1808
    x"D8",x"4C",x"70",x"B7",x"A9",x"00",x"85",x"7D", -- 0x1810
    x"4C",x"AA",x"B7",x"20",x"5B",x"A5",x"A9",x"26", -- 0x1818
    x"85",x"80",x"A9",x"1F",x"85",x"81",x"20",x"A1", -- 0x1820
    x"AC",x"A0",x"03",x"84",x"86",x"B9",x"9D",x"B8", -- 0x1828
    x"99",x"0A",x"90",x"88",x"10",x"F7",x"AD",x"0E", -- 0x1830
    x"90",x"09",x"0F",x"8D",x"0E",x"90",x"A2",x"0F", -- 0x1838
    x"A0",x"90",x"88",x"D0",x"FD",x"C6",x"86",x"D0", -- 0x1840
    x"F7",x"A9",x"0F",x"85",x"86",x"EE",x"0C",x"90", -- 0x1848
    x"88",x"D0",x"FD",x"EA",x"CA",x"D0",x"E9",x"8A", -- 0x1850
    x"8D",x"0C",x"90",x"AD",x"0E",x"90",x"09",x"0F", -- 0x1858
    x"8D",x"0E",x"90",x"20",x"C4",x"B2",x"EA",x"EA", -- 0x1860
    x"C6",x"9F",x"F0",x"0A",x"A4",x"E1",x"B9",x"1E", -- 0x1868
    x"BE",x"30",x"8A",x"4C",x"73",x"B7",x"A2",x"07", -- 0x1870
    x"BD",x"74",x"BB",x"BC",x"93",x"BB",x"99",x"25", -- 0x1878
    x"1F",x"A9",x"00",x"99",x"25",x"97",x"CA",x"10", -- 0x1880
    x"EF",x"20",x"C4",x"B2",x"AD",x"3C",x"18",x"F0", -- 0x1888
    x"03",x"20",x"09",x"A0",x"20",x"C4",x"B2",x"EE", -- 0x1890
    x"3F",x"18",x"4C",x"C3",x"A0",x"00",x"00",x"EF", -- 0x1898
    x"00",x"AE",x"26",x"18",x"B5",x"C0",x"C5",x"90", -- 0x18A0
    x"F0",x"05",x"CA",x"10",x"F7",x"30",x"08",x"B5", -- 0x18A8
    x"D0",x"C5",x"91",x"D0",x"F5",x"F0",x"13",x"A6", -- 0x18B0
    x"7F",x"B5",x"20",x"C5",x"90",x"F0",x"05",x"CA", -- 0x18B8
    x"10",x"F7",x"30",x"08",x"B5",x"28",x"C5",x"91", -- 0x18C0
    x"D0",x"F5",x"E6",x"9D",x"60",x"A4",x"E1",x"BE", -- 0x18C8
    x"2D",x"BE",x"BD",x"FC",x"BF",x"8D",x"00",x"18", -- 0x18D0
    x"BD",x"FE",x"BF",x"8D",x"01",x"18",x"BD",x"E4", -- 0x18D8
    x"BC",x"8D",x"02",x"18",x"BD",x"E6",x"BC",x"8D", -- 0x18E0
    x"03",x"18",x"BD",x"E8",x"BC",x"8D",x"04",x"18", -- 0x18E8
    x"BD",x"EA",x"BC",x"8D",x"05",x"18",x"B9",x"F1", -- 0x18F0
    x"BD",x"85",x"7F",x"B9",x"0F",x"BE",x"8D",x"26", -- 0x18F8
    x"18",x"A9",x"00",x"8D",x"22",x"18",x"A2",x"09", -- 0x1900
    x"8E",x"21",x"18",x"4C",x"F9",x"B2",x"01",x"0D", -- 0x1908
    x"1F",x"1F",x"1F",x"0F",x"03",x"03",x"00",x"60", -- 0x1910
    x"F0",x"F0",x"F0",x"E0",x"80",x"80",x"03",x"07", -- 0x1918
    x"07",x"07",x"03",x"01",x"01",x"00",x"80",x"C0", -- 0x1920
    x"C0",x"C0",x"80",x"00",x"00",x"80",x"00",x"00", -- 0x1928
    x"00",x"00",x"00",x"07",x"0F",x"0F",x"00",x"00", -- 0x1930
    x"00",x"1C",x"3E",x"3E",x"FC",x"FF",x"3F",x"4F", -- 0x1938
    x"07",x"00",x"00",x"00",x"00",x"00",x"FF",x"FC", -- 0x1940
    x"3E",x"3E",x"1C",x"00",x"00",x"00",x"01",x"00", -- 0x1948
    x"00",x"01",x"03",x"03",x"03",x"01",x"00",x"80", -- 0x1950
    x"80",x"C0",x"E0",x"E0",x"E0",x"C0",x"01",x"01", -- 0x1958
    x"07",x"0F",x"0F",x"0F",x"06",x"00",x"C0",x"C0", -- 0x1960
    x"F0",x"F8",x"F8",x"F8",x"B0",x"80",x"00",x"00", -- 0x1968
    x"00",x"38",x"7C",x"7C",x"3F",x"FF",x"00",x"00", -- 0x1970
    x"00",x"00",x"00",x"E0",x"F2",x"FC",x"FF",x"3F", -- 0x1978
    x"7C",x"7C",x"38",x"00",x"00",x"00",x"F0",x"F0", -- 0x1980
    x"E0",x"00",x"00",x"00",x"00",x"00",x"02",x"07", -- 0x1988
    x"0D",x"1F",x"3F",x"5B",x"FF",x"FF",x"00",x"00", -- 0x1990
    x"80",x"C0",x"E0",x"B0",x"F8",x"FC",x"F7",x"9C", -- 0x1998
    x"FE",x"F8",x"DC",x"FE",x"F4",x"FE",x"00",x"00", -- 0x19A0
    x"60",x"95",x"22",x"45",x"F0",x"00",x"00",x"00", -- 0x19A8
    x"10",x"10",x"38",x"FE",x"38",x"10",x"40",x"E0", -- 0x19B0
    x"40",x"00",x"00",x"02",x"07",x"82",x"11",x"40", -- 0x19B8
    x"E0",x"40",x"00",x"08",x"1C",x"08",x"C0",x"90", -- 0x19C0
    x"10",x"38",x"FE",x"38",x"10",x"10",x"04",x"06", -- 0x19C8
    x"07",x"05",x"07",x"07",x"03",x"03",x"20",x"60", -- 0x19D0
    x"E0",x"A0",x"E0",x"E0",x"C0",x"C0",x"07",x"07", -- 0x19D8
    x"07",x"1F",x"1F",x"5F",x"8F",x"7F",x"E0",x"E0", -- 0x19E0
    x"E0",x"F8",x"F8",x"F8",x"F0",x"E0",x"00",x"80", -- 0x19E8
    x"42",x"3B",x"00",x"EE",x"88",x"EE",x"00",x"01", -- 0x19F0
    x"46",x"D8",x"00",x"E9",x"8A",x"EC",x"88",x"EE", -- 0x19F8
    x"00",x"1F",x"24",x"48",x"80",x"00",x"8A",x"E9", -- 0x1A00
    x"00",x"F8",x"24",x"12",x"01",x"00",x"00",x"00", -- 0x1A08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A20
    x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0", -- 0x1A28
    x"F0",x"F0",x"00",x"00",x"00",x"00",x"0F",x"0F", -- 0x1A30
    x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A38
    x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"00",x"00", -- 0x1A40
    x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"F0",x"90", -- 0x1A48
    x"90",x"F0",x"00",x"00",x"00",x"00",x"0F",x"09", -- 0x1A50
    x"09",x"0F",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A58
    x"00",x"00",x"F0",x"90",x"90",x"F0",x"00",x"00", -- 0x1A60
    x"00",x"00",x"0F",x"09",x"09",x"0F",x"90",x"60", -- 0x1A68
    x"60",x"90",x"00",x"00",x"00",x"00",x"09",x"06", -- 0x1A70
    x"06",x"09",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A78
    x"00",x"00",x"90",x"60",x"60",x"90",x"00",x"00", -- 0x1A80
    x"00",x"00",x"09",x"06",x"06",x"09",x"A9",x"FF", -- 0x1A88
    x"8D",x"21",x"91",x"A9",x"01",x"85",x"7D",x"AD", -- 0x1A90
    x"24",x"91",x"AD",x"3F",x"18",x"60",x"AA",x"AA", -- 0x1A98
    x"A9",x"EF",x"8D",x"20",x"91",x"AD",x"21",x"91", -- 0x1AA0
    x"29",x"80",x"F0",x"0A",x"AD",x"1F",x"91",x"CD", -- 0x1AA8
    x"1F",x"91",x"D0",x"F8",x"29",x"20",x"60",x"A9", -- 0x1AB0
    x"FF",x"8D",x"21",x"91",x"A9",x"01",x"85",x"7D", -- 0x1AB8
    x"AD",x"24",x"91",x"AD",x"3F",x"18",x"FF",x"00", -- 0x1AC0
    x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"7F", -- 0x1AC8
    x"7F",x"7F",x"7F",x"7F",x"7F",x"FF",x"FF",x"3F", -- 0x1AD0
    x"3F",x"3F",x"3F",x"3F",x"3F",x"FF",x"FF",x"1F", -- 0x1AD8
    x"1F",x"1F",x"1F",x"1F",x"1F",x"FF",x"FF",x"0F", -- 0x1AE0
    x"0F",x"0F",x"0F",x"0F",x"0F",x"FF",x"FF",x"07", -- 0x1AE8
    x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"03", -- 0x1AF0
    x"03",x"03",x"03",x"03",x"03",x"FF",x"FF",x"01", -- 0x1AF8
    x"01",x"01",x"01",x"01",x"01",x"FF",x"00",x"00", -- 0x1B00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01", -- 0x1B08
    x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09", -- 0x1B10
    x"6E",x"84",x"9A",x"B0",x"C6",x"DC",x"F2",x"08", -- 0x1B18
    x"1E",x"34",x"4A",x"60",x"76",x"8C",x"A2",x"B8", -- 0x1B20
    x"CE",x"E4",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E", -- 0x1B28
    x"1E",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F", -- 0x1B30
    x"1F",x"1F",x"1F",x"1F",x"FD",x"FB",x"EF",x"FB", -- 0x1B38
    x"20",x"40",x"20",x"20",x"04",x"08",x"10",x"00", -- 0x1B40
    x"02",x"03",x"EF",x"7F",x"FB",x"F7",x"80",x"40", -- 0x1B48
    x"20",x"10",x"08",x"04",x"02",x"01",x"93",x"83", -- 0x1B50
    x"8F",x"92",x"85",x"94",x"89",x"8D",x"85",x"77", -- 0x1B58
    x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77", -- 0x1B60
    x"7E",x"8E",x"85",x"98",x"94",x"8D",x"85",x"81", -- 0x1B68
    x"8C",x"92",x"8E",x"84",x"07",x"01",x"0D",x"05", -- 0x1B70
    x"0F",x"16",x"05",x"12",x"20",x"20",x"20",x"20", -- 0x1B78
    x"13",x"10",x"05",x"05",x"04",x"20",x"12",x"15", -- 0x1B80
    x"0E",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x1B88
    x"0E",x"0F",x"2E",x"00",x"01",x"02",x"03",x"16", -- 0x1B90
    x"17",x"18",x"19",x"90",x"95",x"93",x"88",x"A7", -- 0x1B98
    x"86",x"B1",x"A7",x"A0",x"94",x"8F",x"A0",x"92", -- 0x1BA0
    x"95",x"8E",x"A0",x"82",x"8F",x"8E",x"95",x"93", -- 0x1BA8
    x"A0",x"92",x"81",x"94",x"A0",x"A0",x"A0",x"A0", -- 0x1BB0
    x"86",x"8F",x"92",x"A0",x"B2",x"B0",x"B0",x"B0", -- 0x1BB8
    x"B0",x"A0",x"90",x"94",x"93",x"83",x"8F",x"8D", -- 0x1BC0
    x"8D",x"8F",x"84",x"8F",x"92",x"85",x"A0",x"B1", -- 0x1BC8
    x"B9",x"B8",x"B1",x"93",x"94",x"81",x"92",x"A0", -- 0x1BD0
    x"93",x"83",x"92",x"85",x"85",x"8E",x"8D",x"8F", -- 0x1BD8
    x"96",x"85",x"A0",x"92",x"81",x"94",x"A0",x"A0", -- 0x1BE0
    x"A0",x"00",x"01",x"02",x"03",x"04",x"16",x"17", -- 0x1BE8
    x"18",x"19",x"1A",x"1B",x"20",x"20",x"20",x"20", -- 0x1BF0
    x"13",x"15",x"03",x"03",x"05",x"13",x"13",x"21", -- 0x1BF8
    x"21",x"20",x"20",x"20",x"01",x"20",x"0E",x"05", -- 0x1C00
    x"17",x"20",x"08",x"09",x"07",x"08",x"20",x"13", -- 0x1C08
    x"03",x"0F",x"12",x"05",x"20",x"0E",x"0F",x"17", -- 0x1C10
    x"20",x"14",x"12",x"19",x"20",x"06",x"0F",x"12", -- 0x1C18
    x"20",x"14",x"08",x"05",x"20",x"20",x"17",x"0F", -- 0x1C20
    x"12",x"0C",x"04",x"20",x"12",x"05",x"03",x"0F", -- 0x1C28
    x"12",x"04",x"21",x"20",x"20",x"20",x"20",x"20", -- 0x1C30
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x1C38
    x"20",x"20",x"20",x"20",x"00",x"01",x"16",x"17", -- 0x1C40
    x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47", -- 0x1C48
    x"48",x"49",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F", -- 0x1C50
    x"5C",x"5D",x"5E",x"5F",x"10",x"28",x"52",x"25", -- 0x1C58
    x"1F",x"1F",x"1F",x"1F",x"42",x"46",x"4A",x"4E", -- 0x1C60
    x"43",x"47",x"4B",x"4F",x"40",x"44",x"48",x"4C", -- 0x1C68
    x"41",x"45",x"49",x"4D",x"41",x"45",x"49",x"4D", -- 0x1C70
    x"43",x"47",x"4B",x"4F",x"40",x"44",x"48",x"4C", -- 0x1C78
    x"42",x"46",x"4A",x"4E",x"00",x"02",x"00",x"FE", -- 0x1C80
    x"FE",x"00",x"02",x"00",x"1A",x"1E",x"22",x"26", -- 0x1C88
    x"16",x"1E",x"22",x"26",x"68",x"68",x"68",x"68", -- 0x1C90
    x"68",x"06",x"06",x"06",x"01",x"01",x"01",x"01", -- 0x1C98
    x"00",x"01",x"00",x"01",x"16",x"2E",x"02",x"28", -- 0x1CA0
    x"0A",x"30",x"0C",x"3C",x"28",x"22",x"02",x"16", -- 0x1CA8
    x"02",x"0E",x"38",x"0C",x"0C",x"0C",x"1E",x"1E", -- 0x1CB0
    x"20",x"24",x"2A",x"2C",x"2E",x"38",x"3C",x"42", -- 0x1CB8
    x"48",x"56",x"58",x"6A",x"30",x"2C",x"3E",x"0C", -- 0x1CC0
    x"28",x"2A",x"1E",x"2C",x"3E",x"18",x"10",x"26", -- 0x1CC8
    x"34",x"06",x"2E",x"3A",x"06",x"16",x"16",x"1E", -- 0x1CD0
    x"20",x"30",x"3A",x"40",x"40",x"48",x"50",x"50", -- 0x1CD8
    x"50",x"54",x"60",x"64",x"A4",x"C4",x"BC",x"BC", -- 0x1CE0
    x"B4",x"D4",x"BC",x"BC",x"DE",x"E0",x"E3",x"E3", -- 0x1CE8
    x"E0",x"DA",x"D6",x"00",x"ED",x"EF",x"ED",x"00", -- 0x1CF0
    x"EB",x"00",x"EB",x"00",x"F0",x"00",x"EF",x"ED", -- 0x1CF8
    x"EF",x"00",x"F0",x"00",x"F0",x"00",x"EB",x"00", -- 0x1D00
    x"00",x"00",x"00",x"00",x"E0",x"00",x"E3",x"00", -- 0x1D08
    x"E3",x"00",x"E7",x"00",x"E7",x"00",x"EB",x"00", -- 0x1D10
    x"BF",x"CF",x"DD",x"E6",x"E7",x"E8",x"EB",x"ED", -- 0x1D18
    x"BF",x"CF",x"DD",x"E6",x"E7",x"E8",x"EB",x"ED", -- 0x1D20
    x"BF",x"CF",x"DD",x"E6",x"E7",x"E8",x"EB",x"ED", -- 0x1D28
    x"BF",x"CF",x"DD",x"E6",x"E7",x"E8",x"EB",x"ED", -- 0x1D30
    x"00",x"DC",x"DA",x"D8",x"D6",x"DE",x"DC",x"DA", -- 0x1D38
    x"D8",x"D6",x"DE",x"DC",x"DA",x"D8",x"D6",x"D5", -- 0x1D40
    x"00",x"00",x"00",x"00",x"CE",x"D0",x"00",x"D0", -- 0x1D48
    x"00",x"00",x"D6",x"00",x"00",x"00",x"00",x"00", -- 0x1D50
    x"CE",x"D0",x"00",x"D0",x"00",x"00",x"D6",x"00", -- 0x1D58
    x"00",x"00",x"00",x"00",x"C0",x"00",x"00",x"C8", -- 0x1D60
    x"00",x"00",x"CE",x"00",x"00",x"00",x"00",x"00", -- 0x1D68
    x"C0",x"00",x"00",x"C8",x"00",x"00",x"CE",x"00", -- 0x1D70
    x"DB",x"00",x"DB",x"DF",x"E7",x"E4",x"E3",x"E7", -- 0x1D78
    x"E3",x"EA",x"EC",x"ED",x"EF",x"D5",x"00",x"D5", -- 0x1D80
    x"DB",x"E4",x"E7",x"E3",x"ED",x"E3",x"E7",x"DB", -- 0x1D88
    x"00",x"E7",x"E1",x"E7",x"E3",x"EA",x"EC",x"E4", -- 0x1D90
    x"DF",x"E4",x"00",x"E4",x"E7",x"E4",x"E7",x"E3", -- 0x1D98
    x"ED",x"E3",x"E7",x"E3",x"01",x"02",x"01",x"02", -- 0x1DA0
    x"01",x"02",x"01",x"02",x"01",x"02",x"01",x"02", -- 0x1DA8
    x"01",x"02",x"03",x"04",x"02",x"01",x"05",x"01", -- 0x1DB0
    x"02",x"03",x"01",x"02",x"03",x"04",x"02",x"01", -- 0x1DB8
    x"05",x"01",x"02",x"03",x"01",x"02",x"03",x"04", -- 0x1DC0
    x"02",x"01",x"05",x"01",x"02",x"03",x"01",x"02", -- 0x1DC8
    x"03",x"DB",x"DB",x"CF",x"DF",x"DB",x"E7",x"EA", -- 0x1DD0
    x"ED",x"E4",x"ED",x"E4",x"ED",x"DB",x"E7",x"DB", -- 0x1DD8
    x"DB",x"CF",x"E7",x"E3",x"DB",x"DF",x"E7",x"DF", -- 0x1DE0
    x"E7",x"D9",x"E7",x"D9",x"E7",x"D9",x"E7",x"DB", -- 0x1DE8
    x"E7",x"02",x"03",x"06",x"03",x"04",x"05",x"07", -- 0x1DF0
    x"04",x"05",x"06",x"06",x"06",x"06",x"07",x"07", -- 0x1DF8
    x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"05", -- 0x1E00
    x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"07", -- 0x1E08
    x"07",x"0F",x"07",x"07",x"07",x"0F",x"07",x"07", -- 0x1E10
    x"07",x"0F",x"07",x"07",x"07",x"0F",x"00",x"00", -- 0x1E18
    x"FF",x"00",x"00",x"00",x"FF",x"00",x"00",x"00", -- 0x1E20
    x"FF",x"00",x"00",x"00",x"FF",x"00",x"00",x"00", -- 0x1E28
    x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00", -- 0x1E30
    x"01",x"01",x"01",x"01",x"00",x"0F",x"F0",x"00", -- 0x1E38
    x"7F",x"CC",x"33",x"FA",x"40",x"4D",x"B3",x"FA", -- 0x1E40
    x"5B",x"41",x"80",x"02",x"11",x"0D",x"E1",x"F2", -- 0x1E48
    x"11",x"0D",x"E9",x"82",x"5B",x"41",x"88",x"1A", -- 0x1E50
    x"40",x"4D",x"B8",x"C0",x"7F",x"CC",x"38",x"1E", -- 0x1E58
    x"00",x"0C",x"00",x"FE",x"3C",x"0C",x"7C",x"00", -- 0x1E60
    x"20",x"C0",x"00",x"00",x"2E",x"DA",x"DD",x"BE", -- 0x1E68
    x"2E",x"DA",x"DD",x"3E",x"20",x"C2",x"9D",x"06", -- 0x1E70
    x"28",x"02",x"01",x"06",x"0B",x"3E",x"D1",x"B6", -- 0x1E78
    x"BA",x"00",x"D4",x"30",x"9A",x"F4",x"D4",x"3E", -- 0x1E80
    x"9A",x"C4",x"17",x"BE",x"82",x"04",x"17",x"80", -- 0x1E88
    x"82",x"C4",x"90",x"00",x"92",x"F4",x"97",x"21", -- 0x1E90
    x"90",x"04",x"90",x"21",x"90",x"E4",x"D6",x"AD", -- 0x1E98
    x"1E",x"E0",x"56",x"AD",x"00",x"E7",x"56",x"A1", -- 0x1EA0
    x"4E",x"E7",x"40",x"A1",x"4E",x"E0",x"1F",x"AD", -- 0x1EA8
    x"40",x"02",x"40",x"2D",x"70",x"3A",x"47",x"A1", -- 0x1EB0
    x"73",x"80",x"07",x"A1",x"73",x"FC",x"00",x"00", -- 0x1EB8
    x"40",x"0C",x"F1",x"EC",x"5A",x"00",x"80",x"2C", -- 0x1EC0
    x"5A",x"9E",x"8E",x"2C",x"1A",x"80",x"A0",x"A0", -- 0x1EC8
    x"42",x"9E",x"A0",x"AC",x"5E",x"9E",x"8E",x"2C", -- 0x1ED0
    x"50",x"80",x"80",x"2C",x"50",x"B8",x"F1",x"EC", -- 0x1ED8
    x"57",x"B8",x"00",x"00",x"47",x"80",x"FC",x"9C", -- 0x1EE0
    x"70",x"00",x"00",x"9C",x"71",x"A0",x"0B",x"80", -- 0x1EE8
    x"71",x"AA",x"AB",x"BE",x"00",x"2A",x"A8",x"3E", -- 0x1EF0
    x"61",x"AA",x"AB",x"06",x"6F",x"AA",x"AB",x"36", -- 0x1EF8
    x"00",x"00",x"00",x"00",x"DD",x"AA",x"AB",x"00", -- 0x1F00
    x"DD",x"AA",x"AB",x"3E",x"0C",x"2A",x"A8",x"3E", -- 0x1F08
    x"61",x"AA",x"AB",x"06",x"6F",x"A0",x"0B",x"36", -- 0x1F10
    x"00",x"00",x"00",x"00",x"00",x"0F",x"F0",x"00", -- 0x1F18
    x"7F",x"CC",x"33",x"FA",x"40",x"4D",x"B3",x"FA", -- 0x1F20
    x"5B",x"41",x"80",x"02",x"11",x"07",x"E1",x"F2", -- 0x1F28
    x"11",x"07",x"E9",x"82",x"5B",x"41",x"88",x"1A", -- 0x1F30
    x"40",x"4D",x"B8",x"C0",x"7F",x"CC",x"38",x"1E", -- 0x1F38
    x"00",x"0C",x"00",x"FE",x"3C",x"0C",x"7C",x"00", -- 0x1F40
    x"20",x"C0",x"00",x"00",x"27",x"FA",x"DD",x"BE", -- 0x1F48
    x"27",x"FA",x"DD",x"3E",x"20",x"C2",x"9D",x"06", -- 0x1F50
    x"28",x"02",x"01",x"06",x"0B",x"3E",x"D1",x"B6", -- 0x1F58
    x"BA",x"00",x"D4",x"30",x"9A",x"F4",x"D4",x"3E", -- 0x1F60
    x"9A",x"C4",x"17",x"BE",x"82",x"14",x"17",x"80", -- 0x1F68
    x"82",x"C4",x"90",x"00",x"92",x"F4",x"9F",x"21", -- 0x1F70
    x"90",x"04",x"90",x"2D",x"90",x"E4",x"D6",x"AD", -- 0x1F78
    x"1E",x"80",x"56",x"A1",x"00",x"8F",x"56",x"BF", -- 0x1F80
    x"4E",x"EF",x"40",x"BF",x"4E",x"E0",x"1F",x"A1", -- 0x1F88
    x"40",x"22",x"40",x"2D",x"70",x"3A",x"47",x"AD", -- 0x1F90
    x"73",x"80",x"07",x"A1",x"73",x"FC",x"00",x"00", -- 0x1F98
    x"40",x"0C",x"FD",x"EC",x"5A",x"00",x"80",x"2C", -- 0x1FA0
    x"5A",x"FE",x"AE",x"AC",x"1A",x"80",x"A0",x"A0", -- 0x1FA8
    x"42",x"9E",x"A0",x"AC",x"5E",x"9E",x"BE",x"AC", -- 0x1FB0
    x"50",x"80",x"80",x"2C",x"50",x"B8",x"F7",x"EC", -- 0x1FB8
    x"57",x"B8",x"00",x"00",x"47",x"80",x"FC",x"9C", -- 0x1FC0
    x"70",x"00",x"00",x"9C",x"71",x"AA",x"AB",x"80", -- 0x1FC8
    x"71",x"AA",x"AB",x"BE",x"00",x"2A",x"A8",x"3E", -- 0x1FD0
    x"61",x"AA",x"AB",x"06",x"6F",x"AA",x"AB",x"36", -- 0x1FD8
    x"00",x"00",x"00",x"00",x"DD",x"AA",x"AB",x"00", -- 0x1FE0
    x"DD",x"AA",x"AB",x"3E",x"0C",x"2A",x"A8",x"3E", -- 0x1FE8
    x"61",x"AA",x"AB",x"06",x"6F",x"AA",x"AB",x"36", -- 0x1FF0
    x"00",x"00",x"00",x"00",x"3C",x"1C",x"BE",x"BF"  -- 0x1FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
